* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param GAU = AGAUSS(0,0.05537,1)
.param GAU2 = AGAUSS(0,0.01662,1)
.param sky130_fd_pr__pnp_05v5_W0p68L0p68__bf_slope = 0.0
.param sky130_fd_pr__pnp_05v5_W0p68L0p68__is_slope = 0.0
* statistics '
*   mismatch '
*     vary  sky130_fd_pr__pnp_05v5_W0p68L0p68__bf_slope dist=gauss std=0.05537
*     vary  sky130_fd_pr__pnp_05v5_W0p68L0p68__is_slope dist=gauss std=0.01662
*   '
* '
.subckt  sky130_fd_pr__pnp_05v5_W0p68L0p68 Collector Base Emitter
+ 
.param  mult = 1.0
*(mismatch parameter sky130_fd_pr__pnp_05v5_W0p68L0p68__bf_slope)
+ sky130_fd_pr__pnp_05v5_W0p68L0p68__bf_mm = '(19.35*dkbfpp*MC_MM_SWITCH*GAU/sqrt(mult))'
*(mismatch parameter sky130_fd_pr__pnp_05v5_W0p68L0p68__is_slope)
+ sky130_fd_pr__pnp_05v5_W0p68L0p68__is_mm = '(1.5075e-018*dkispp*MC_MM_SWITCH*GAU2/sqrt(mult))'
qsky130_fd_pr__pnp_05v5_W0p68L0p68 Collector Base Emitter Collector sky130_fd_pr__pnp_05v5_W0p68L0p68__model
.model sky130_fd_pr__pnp_05v5_W0p68L0p68__model pnp level = 1.0
* General Parameters
+ tref = 30.0
* Capacitance Parameters
+ cjc = 6.255e-015 cje = 6.113e-016 cjs = 0.0
+ fc = 0.5 mjc = 0.24 mje = 0.3 mjs = 0.24
+ vjc = 0.54 vje = 0.74 vjs = 0.54 xcjc = 1.0
+ ptf = 0 tf = 6.15385e-010 tr = 5e-008 vtf = 1.0e-12
+ xtf = 0.0
* Noise Parameters
+ af = 1.60722 kf = 4.9435066e-11
* DC Parameters
+ is = '1.5075e-018*1.00*dkispp+sky130_fd_pr__pnp_05v5_W0p68L0p68__is_mm' rb = 316.21 re = 219 irb = 0.027411
+ rc = 531 rbm = 243.58 bf = '19.35*dkbfpp+sky130_fd_pr__pnp_05v5_W0p68L0p68__bf_mm' nf = '1.028*dknfpp'
+ vaf = 152.06 ikf = 3.3057e-005 ise = 9.4936e-017 ne = 1.6444
+ ns = 1 br = 0.2675 iss = 0 nr = 1.0
+ var = 4.3 ikr = 0.00043 nkf = 0.5 isc = 1.2e-15
+ nc = 1.003
* Temperature Parameters
+ xtb = 2.2132 xti = 1.1 eg = 1.2 tikf1 = -0.0037823
+ tnf1 = 1.972e-006 tnf2 = -8.8e-7
.ends sky130_fd_pr__pnp_05v5_W0p68L0p68
