* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param GAU = AGAUSS(0,1.0,1)
.param npnpolyhv_is_slope_spectre = 0.0
.param npnpolyhv_bf_slope_spectre = 0.0
* statistics {
*   mismatch {
*     vary  npnpolyhv_is_slope_spectre dist=gauss std=1.0
*     vary  npnpolyhv_bf_slope_spectre dist=gauss std=1.0
*   }
* }
.subckt  sky130_fd_pr__npn_11v0_W1p00L1p00 c b e s
+ 
.param  mult = 1.0
qsky130_fd_pr__npn_11v0_W1p00L1p00 c1 b e s sky130_fd_pr__npn_11v0_W1p00L1p00__base
rc c c1 r = 440 tc1 = -4.0e-3
q2 s c1 b s sky130_fd_pr__pnp_05v5_W0p68L0p68__polyhv
d1 s b sky130_fd_pr__model__parasitic__diode_ps2dn area = 1.34
.model sky130_fd_pr__npn_11v0_W1p00L1p00__base npn level = 1.0
* General Parameters
+ tref = 30.0
* Capacitance Parameters
+ dcap = 2 cjc = '1.60339e-014*sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult' cje = '10.30981e-015*sky130_fd_pr__nfet_01v8__ajunction_mult'
+ cjs = '3.05951e-014*sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult' fc = 0.5 mjc = 0.33982 mje = 0.44
+ mjs = 0.49 vjc = 0.58758 vje = 0.729 vjs = 0.5348
+ xcjc = 1 itf = 9.6e-03 ptf = 20 tf = 10.84e-11
+ tr = 0 vtf = 0.5 xtf = 2.9
* Noise Parameters
+ af = 1.9 kf = 5.0e-10
* DC Parameters
*(mismatch parameter npnpolyhv_is_slope_spectre)
+ is = '1.1082e-017*dkisnpnpolyhv + 1.1082e-017*dkisnpnpolyhv*0.003/sqrt(mult)*MC_MM_SWITCH*GAU' rb = 1400.0
+ re = 85 irb = 4.424e-005 rc = 1.0 rbm = 400.07
*(mismatch parameter npnpolyhv_bf_slope_spectre)
+ bf = '141.286*dkbfnpnpolyhv + 141.286*dkbfnpnpolyhv*0.05/sqrt(mult)*MC_MM_SWITCH*GAU' nf = 1.0262306 vaf = 100 ikf = 0.00046731
+ ise = 5.3935e-016 ne = 1.7527 ns = 1 br = 100.0
+ iss = 0 nr = 1.0262306
+ var = 0 ikr = 0.00046731 nkf = 0.31875 isc = 0.0
+ nc = 2.0
* Temperature Parameters
+ xtb = 0 xti = 2.7498 eg = 1.1714 gap1 = 0.0
+ gap2 = 0 ctc = 0 cte = 0 cts = 0.0
+ tlev = 0 tlevc = 0 tvjc = 0 tvje = 0.0
+ tvjs = 0 tis1 = 0 tise1 = 0 tisc1 = 0.0
+ tnf1 = 4.208e-005 tnr1 = -0.000522 tne1 = 0 tnc1 = 0.0
+ tbf1 = 7.4942e-003 tbr1 = 0 tiss1 = 0 tvaf1 = 0.0
+ tvar1 = 0 tikf1 = -0.012219846 tikr1 = 0 tns1 = 0.0
+ trb1 = -0.0029419354 trc1 = 3.7260032e-005 tre1 = 5e-3 tirb1 = 0.0
+ trm1 = 0.004459028 tmjc1 = 0 tmje1 = 0 tmjs1 = 0.0
+ ttf1 = 0 titf1 = 0 ttr1 = 0 tis2 = 4.0e-12
+ tise2 = 0 tisc2 = 0 tnf2 = -3.372e-007 tnr2 = 1.8e-6
+ tne2 = 0 tnc2 = 0 tbf2 = 7.633e-006 tbr2 = 0.0
+ tiss2 = 0 tvaf2 = 0 tvar2 = 0 tikf2 = 9.3646292e-5
+ tikr2 = 0 tns2 = 0 trb2 = 3.4143764e-005 trc2 = 3.0650517e-7
+ tre2 = 0.0 tirb2 = 0 trm2 = -4.9458296e-005 tmjc2 = 0.0
+ tmje2 = 0 tmjs2 = 0 ttf2 = 0 titf2 = 0.0
+ ttr2 = 0.0
.model sky130_fd_pr__pnp_05v5_W0p68L0p68__polyhv pnp level = 1.0
* General Parameters
+ tref = 30.0
* Capacitance Parameters
+ dcap = 2 cjc = 0 cje = 0.0
+ cjs = 0 fc = 0.5 mjc = 0.33 mje = 0.33
+ mjs = 0.5 vjc = 0.75 vje = 0.75 vjs = 0.75
+ xcjc = 1.0
+ itf = 0 ptf = 0 tf = 0 tr = 0.0
+ vtf = 0.5 xtf = 0.0
* Noise Parameters
+ af = 1.9 kf = 5.0e-9
* DC Parameters
*(mismatch parameter npnpolyhv_is_slope_spectre)
+ is = '1.2252871e-016*dkisnpnpolyhv + 1.2252871e-016*dkisnpnpolyhv*0.003/sqrt(mult)*MC_MM_SWITCH*GAU' rb = 1922.4
+ re = 6000 irb = 0 rc = 1 rbm = 46.144
*(mismatch parameter npnpolyhv_bf_slope_spectre)
+ bf = '25*dkbfnpnpolyhv + 25*dkbfnpnpolyhv*0.05/sqrt(mult)*MC_MM_SWITCH*GAU' nf = 1.0161516 vaf = 0 ikf = 100.0
+ ise = 1e-016 ne = 2 ns = 1 br = 1.0
+ ibc = 0 iss = 0 nr = 1.0
+ var = 0 ikr = 1e-10 nkf = 0.41826 isc = 0.0
+ nc = 2.0
* Temperature Parameters
+ xtb = 0 xti = 5.351377 eg = 1.11 gap1 = 0.0
+ gap2 = 0 ctc = 0.0
+ cte = 0 cts = 0 tlev = 0 tlevc = 0.0
+ tvjc = 0 tvje = 0 tvjs = 0.0
+ tis1 = 0 tise1 = 0 tisc1 = 0.0
+ tnf1 = -6e-3 tnr1 = 0 tne1 = 0 tnc1 = 0.0
+ tbf1 = 0 tbr1 = 0 tiss1 = 0 tvaf1 = 0.0
+ tvar1 = 0 tikf1 = 0 tikr1 = 0 tns1 = 0.0
+ trb1 = 0 trc1 = 0 tre1 = -0.005 tirb1 = 0.0
+ trm1 = 0 tmjc1 = 0 tmje1 = 0 tmjs1 = 0.0
+ ttf1 = 0 titf1 = 0 ttr1 = 0 tis2 = 0.0
+ tise2 = 0 tisc2 = 0 tnf2 = 0 tnr2 = 0.0
+ tne2 = 0 tnc2 = 0 tbf2 = 0 tbr2 = 0.0
+ tiss2 = 0 tvaf2 = 0 tvar2 = 0 tikf2 = 0.0
+ tikr2 = 0 tns2 = 0 trb2 = 0 trc2 = 0.0
+ tre2 = 0 tirb2 = 0 trm2 = 0 tmjc2 = 0.0
+ tmje2 = 0 tmjs2 = 0 ttf2 = 0 titf2 = 0.0
+ ttr2 = 0.0
.ends sky130_fd_pr__npn_11v0_W1p00L1p00
