* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param GAU = AGAUSS(0,1.0,1)
.param
+ sky130_fd_pr__pfet_g5v0d16v0__mm_mult = 0.9
.param sky130_fd_pr__pfet_g5v0d16v0__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d16v0__wint_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d16v0__lint_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d16v0__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d16v0__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d16v0__nfactor_slope_spectre = 0.0
* statistics '
*   process '
*   '
*   mismatch '
*     vary sky130_fd_pr__pfet_g5v0d16v0__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d16v0__wint_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d16v0__lint_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d16v0__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d16v0__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d16v0__nfactor_slope_spectre dist=gauss std = 1.0
*   '
* '
.subckt  sky130_fd_pr__pfet_g5v0d16v0__base d g s b
+ 
.param  l = 1 w = 1 nf = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 delvto = 0.0
msky130_fd_pr__pfet_g5v0d16v0__base d g s b sky130_fd_pr__pfet_g5v0d16v0__model_base l = 'l' w = 'w' nf = 'nf' ad = 'ad' as = 'as' pd = 'pd' ps = 'ps' nrd = 'nrd' nrs = 'nrs' sa = 'sa' sb = 'sb' sd = 'sd'
.model sky130_fd_pr__pfet_g5v0d16v0__model_base.0 pmos
* Model Flag Parameters
+ lmin = 0.655e-06 lmax = 0.665e-06 wmin = 4.990000e-006 wmax = 5.010000e-5
+ level = 5.400000e+1
+ version = 4.500000e+0
+ binunit = 2.000000e+0
+ mobmod = .000000e+0
+ capmod = 2.000000e+0
+ igcmod = .000000e+0
+ igbmod = .000000e+0
+ geomod = .000000e+0
+ diomod = 1.000000e+0
+ rdsmod = 1.000000e+0
+ rbodymod = 1.000000e+0
+ rgatemod = .000000e+0
+ permod = 1.000000e+0
+ acnqsmod = .000000e+0
+ trnqsmod = .000000e+0
+ fnoimod = 1.000000e+0
+ tnoimod = 1.000000e+0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d16v0__toxe_slope_spectre)
+ toxe = '1.160000e-008*sky130_fd_pr__pfet_g5v0d16v0__toxe_mult+MC_MM_SWITCH*GAU*(1.16e-008*sky130_fd_pr__pfet_g5v0d16v0__toxe_mult*(sky130_fd_pr__pfet_g5v0d16v0__mm_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1+0.05e-2)/sqrt(l*w*mult)))'
+ toxm = 1.160000e-8
+ epsrox = 3.900000e+0
+ xj = 1.500000e-7
+ ngate = 1.000000e+23
+ ndep = 1.700000e+17
+ nsd = 1.000000e+20
+ rsh = '1.000000e+000*sky130_fd_pr__pfet_g5v0d16v0__rshp_mult'
+ rshg = 1.000000e-1
* Basic Model Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d16v0__wint_slope_spectre)
+ wint = '0.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__wint_diff+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d16v0__mm_mult*sky130_fd_pr__pfet_g5v0d10v5__wint_slope/sqrt(l))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d16v0__lint_slope_spectre)
+ lint = '3.445300e-008+sky130_fd_pr__pfet_g5v0d16v0__lint_diff+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d16v0__mm_mult*sky130_fd_pr__pfet_g5v0d10v5__lint_slope/sqrt(w))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d16v0__vth0_slope_spectre)
+ vth0 = '-1.043500e+000+sky130_fd_pr__pfet_g5v0d16v0__vth0_diff_0+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d16v0__mm_mult*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope+0.0065)/sqrt(l*w*mult))'
+ k1 = 6.831000e-1
+ k2 = '-1.303200e-003+sky130_fd_pr__pfet_g5v0d16v0__k2_diff_0'
+ k3 = .000000e+0
+ k3b = .000000e+0
+ w0 = .000000e+0
+ dvt0 = .000000e+0
+ dvt1 = 5.300000e-1
+ dvt2 = -3.200000e-2
+ dvt0w = .000000e+0
+ dvt1w = 5.300000e+6
+ dvt2w = -3.200000e-2
+ dsub = '3.416000e-001+sky130_fd_pr__pfet_g5v0d16v0__dsub_diff_0'
+ minv = .000000e+0
+ voffl = .000000e+0
+ dvtp0 = .000000e+0
+ dvtp1 = .000000e+0
+ lpe0 = '1.400000e-007+sky130_fd_pr__pfet_g5v0d16v0__lpe0_diff_0'
+ lpeb = -6.500000e-8
+ vbm = -3.000000e+0
+ phin = .000000e+0
+ cdsc = 2.520000e-4
+ cdscb = .000000e+0
+ cdscd = .000000e+0
+ cit = .000000e+0
*(mismatch parameter sky130_fd_pr__pfet_g5v0d16v0__voff_slope_spectre)
+ voff = '-1.372000e-001+sky130_fd_pr__pfet_g5v0d16v0__voff_diff_0+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d16v0__mm_mult*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope+0.02)/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d16v0__nfactor_slope_spectre)
+ nfactor = '7.100000e-001+sky130_fd_pr__pfet_g5v0d16v0__nfactor_diff_0+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d16v0__mm_mult*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope+0.3)/sqrt(l*w*mult))'
+ eta0 = '8.729800e-002+sky130_fd_pr__pfet_g5v0d16v0__eta0_diff_0'
+ etab = -5.000000e-2
+ u0 = '2.707600e-002+sky130_fd_pr__pfet_g5v0d16v0__u0_diff_0'
+ ua = '2.585600e-009+sky130_fd_pr__pfet_g5v0d16v0__ua_diff_0'
+ ub = '4.595800e-019+sky130_fd_pr__pfet_g5v0d16v0__ub_diff_0'
+ uc = -1.220000e-10
+ eu = 1.670000e+0
+ vsat = '7.660800e+004+sky130_fd_pr__pfet_g5v0d16v0__vsat_diff_0'
+ a0 = '3.820000e-001+sky130_fd_pr__pfet_g5v0d16v0__a0_diff_0'
+ ags = '1.291200e-001+sky130_fd_pr__pfet_g5v0d16v0__ags_diff_0'
+ a1 = .000000e+0
+ a2 = 7.200000e-1
+ b0 = '4.000000e-012+sky130_fd_pr__pfet_g5v0d16v0__b0_diff_0'
+ b1 = '0.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__b1_diff_0'
+ keta = '-3.321800e-002+sky130_fd_pr__pfet_g5v0d16v0__keta_diff_0'
+ dwg = .000000e+0
+ dwb = .000000e+0
+ pclm = '1.000000e-001+sky130_fd_pr__pfet_g5v0d16v0__pclm_diff_0'
+ pdiblc1 = 3.900000e-1
+ pdiblc2 = 8.600000e-3
+ pdiblcb = -5.400000e-5
+ drout = 5.600000e-1
+ pvag = 5.040000e-1
+ delta = 8.900000e-3
+ pscbe1 = 5.088000e+8
+ pscbe2 = 6.945200e-9
+ fprout = .000000e+0
+ pdits = '0.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__pdits_diff_0'
+ pditsd = '0.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__pditsd_diff_0'
+ pditsl = .000000e+0
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = '3.310200e+002+sky130_fd_pr__pfet_g5v0d16v0__rdsw_diff_0'
+ rsw = 1.000000e+2
+ rdw = '1.000000e+001+sky130_fd_pr__pfet_g5v0d16v0__rdw_diff_0'
+ rdswmin = .000000e+0
+ rdwmin = .000000e+0
+ rswmin = .000000e+0
+ prwg = .000000e+0
+ prwb = -4.000000e-4
+ wr = 1.000000e+0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.000000e-7
+ alpha1 = 1.001000e+0
+ beta0 = 1.000000e+2
* Gidl Induced Drain Leakage Model Parameters
+ agidl = '1.650000e-010+sky130_fd_pr__pfet_g5v0d16v0__agidl_diff_0'
+ bgidl = '5.999300e+009+sky130_fd_pr__pfet_g5v0d16v0__bgidl_diff_0'
+ cgidl = '1.394000e+000+sky130_fd_pr__pfet_g5v0d16v0__cgidl_diff_0'
+ egidl = 4.920000e-2
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 1.160000e-8
+ aigbacc = '4.300000e-001+sky130_fd_pr__pfet_g5v0d16v0__aigbacc_diff_0'
+ bigbacc = 5.400000e-2
+ cigbacc = 7.500000e-2
+ nigbacc = '1.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__nigbacc_diff_0'
+ aigbinv = '3.500000e-001+sky130_fd_pr__pfet_g5v0d16v0__aigbinv_diff_0'
+ bigbinv = 3.000000e-2
+ cigbinv = 6.000000e-3
+ eigbinv = 1.100000e+0
+ nigbinv = '3.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__nigbinv_diff_0'
+ aigc = '4.300000e-001+sky130_fd_pr__pfet_g5v0d16v0__aigc_diff_0'
+ bigc = 5.400000e-2
+ cigc = 7.500000e-2
+ aigsd = '4.300000e-001+sky130_fd_pr__pfet_g5v0d16v0__aigsd_diff_0'
+ bigsd = '5.400000e-002+sky130_fd_pr__pfet_g5v0d16v0__bigsd_diff_0'
+ cigsd = 7.500000e-2
+ nigc = 1.000000e+0
+ poxedge = 1.000000e+0
+ pigcd = 1.000000e+0
+ ntox = 1.000000e+0
* Charge AND Capacitance Model Parameters
+ dlc = '-9.682600e-008+sky130_fd_pr__pfet_g5v0d16v0__dlc_diff+sky130_fd_pr__pfet_g5v0d16v0__dlc_rotweak'
+ dwc = '0.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__dwc_diff'
+ xpart = .000000e+0
+ cgso = '1.977100e-010*sky130_fd_pr__pfet_g5v0d16v0__soverlap_mult'
+ cgdo = '1.977100e-010*sky130_fd_pr__pfet_g5v0d16v0__doverlap_mult'
+ cgbo = .000000e+0
+ cgdl = '1.117200e-012*sky130_fd_pr__pfet_g5v0d16v0__doverlap_mult'
+ cgsl = '1.152000e-012*sky130_fd_pr__pfet_g5v0d16v0__soverlap_mult'
+ clc = 6.324000e-9
+ cle = 8.910000e-1
+ cf = '0.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__cf_diff'
+ ckappas = 6.000000e-1
+ ckappad = 6.000000e-1
+ vfbcv = -1.000000e+0
+ acde = 9.129800e-1
+ moin = 1.556200e+1
+ noff = 1.045000e+0
+ voffcv = -1.815100e-1
* High-Speed/RF Model Parameters
* Flicker AND Thermal Noise Model Parameters
+ ef = 1.000000e+0
+ noia = 6.250000e+41
+ noib = 3.125000e+26
+ noic = 8.750000e+9
+ em = 4.100000e+7
* Layout-Dependent Parasitics Model Parameters
+ xl = .000000e+0
+ xw = .000000e+0
+ dmcg = .000000e+0
+ dmdg = .000000e+0
+ dmcgt = .000000e+0
+ xgw = .000000e+0
+ xgl = .000000e+0
+ ngcon = 1.000000e+0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.148300e-5
+ jsws = 4.020000e-12
+ jtssws = '4.020000e-012+sky130_fd_pr__pfet_g5v0d16v0__jtssws_diff_0'
+ ijthsfwd = 1.000000e-1
+ ijthsrev = 1.000000e-1
+ bvs = 1.269000e+1
+ xjbvs = 1.000000e+0
+ pbs = 6.587000e-1
+ cjs = '7.754700e-004*sky130_fd_pr__pfet_g5v0d16v0__ajunction_mult'
+ mjs = 3.395600e-1
+ pbsws = 1.000000e+0
+ cjsws = '9.871700e-011*sky130_fd_pr__pfet_g5v0d16v0__pjunction_mult'
+ mjsws = 2.467600e-1
+ pbswgs = 3.000000e+0
+ cjswgs = '1.460000e-010*sky130_fd_pr__pfet_g5v0d16v0__pjunction_mult'
+ mjswgs = 8.100000e-1
* Temperature Dependence Parameters
+ tnom = 3.000000e+1
+ kt1 = '-4.930800e-001+sky130_fd_pr__pfet_g5v0d16v0__kt1_diff_0'
+ kt1l = 1.000000e-11
+ kt2 = 5.633800e-4
+ ute = -1.646200e+0
+ ua1 = 1.218100e-9
+ ub1 = -1.241200e-18
+ uc1 = 8.272000e-12
+ prt = .000000e+0
+ at = -6.400000e+4
+ tvoff = '1.500000e-002+sky130_fd_pr__pfet_g5v0d16v0__tvoff_diff_0'
+ njs = 1.363200e+0
+ njd = 1.079100e+0
+ tpb = 1.671000e-3
+ tcj = 9.600000e-4
+ tpbsw = .000000e+0
+ tcjsw = 3.000000e-5
+ tpbswg = .000000e+0
+ tcjswg = .000000e+0
+ xtis = 1.000000e+1
+ xtid = 3.000000e+0
* DW AND DL Parameters
+ ll = .000000e+0
+ wl = .000000e+0
+ lln = 1.000000e+0
+ wln = 1.000000e+0
+ lw = .000000e+0
+ ww = .000000e+0
+ lwn = 1.000000e+0
+ wwn = 1.000000e+0
+ lwl = .000000e+0
+ wwl = .000000e+0
+ llc = .000000e+0
+ wlc = .000000e+0
+ lwc = .000000e+0
+ wwc = .000000e+0
+ lwlc = .000000e+0
+ wwlc = .000000e+0
* Stress Parameters
+ saref = .28e-6
+ sbref = 1.19e-6
+ kvth0 = '0.0+sky130_fd_pr__pfet_g5v0d16v0__kvth0_diff'
+ lkvth0 = '0.0+sky130_fd_pr__pfet_g5v0d16v0__lkvth0_diff'
+ wkvth0 = '0.0+sky130_fd_pr__pfet_g5v0d16v0__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 1.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0.0+sky130_fd_pr__pfet_g5v0d16v0__ku0_diff'
+ lku0 = '0.0+sky130_fd_pr__pfet_g5v0d16v0__lku0_diff'
+ wku0 = '0.0+sky130_fd_pr__pfet_g5v0d16v0__wku0_diff'
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 1.0
+ wlodku0 = 1.0
+ kvsat = '0.0+sky130_fd_pr__pfet_g5v0d16v0__kvsat_diff'
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_g5v0d16v0__model_base.1 pmos
* Model Flag Parameters
+ lmin = 2.15e-06 lmax = 2.17e-06 wmin = 4.990000e-006 wmax = 5.010000e-5
+ level = 5.400000e+1
+ version = 4.500000e+0
+ binunit = 2.000000e+0
+ mobmod = .000000e+0
+ capmod = 2.000000e+0
+ igcmod = .000000e+0
+ igbmod = .000000e+0
+ geomod = .000000e+0
+ diomod = 1.000000e+0
+ rdsmod = 1.000000e+0
+ rbodymod = 1.000000e+0
+ rgatemod = .000000e+0
+ permod = 1.000000e+0
+ acnqsmod = .000000e+0
+ trnqsmod = .000000e+0
+ fnoimod = 1.000000e+0
+ tnoimod = 1.000000e+0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d16v0__toxe_slope_spectre)
+ toxe = '1.160000e-008*sky130_fd_pr__pfet_g5v0d16v0__toxe_mult+MC_MM_SWITCH*GAU*(1.16e-008*sky130_fd_pr__pfet_g5v0d16v0__toxe_mult*(sky130_fd_pr__pfet_g5v0d16v0__mm_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope2+0.03e-2)/sqrt(l*w*mult)))'
+ toxm = 1.160000e-8
+ epsrox = 3.900000e+0
+ xj = 1.500000e-7
+ ngate = 1.000000e+23
+ ndep = 1.700000e+17
+ nsd = 1.000000e+20
+ rsh = '1.000000e+000*sky130_fd_pr__pfet_g5v0d16v0__rshp_mult'
+ rshg = 1.000000e-1
* Basic Model Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d16v0__wint_slope_spectre)
+ wint = '0.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__wint_diff+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d16v0__mm_mult*sky130_fd_pr__pfet_g5v0d10v5__wint_slope/sqrt(l))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d16v0__lint_slope_spectre)
+ lint = '3.445300e-008+sky130_fd_pr__pfet_g5v0d16v0__lint_diff+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d16v0__mm_mult*sky130_fd_pr__pfet_g5v0d10v5__lint_slope/sqrt(w))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d16v0__vth0_slope_spectre)
+ vth0 = '-1.043500e+000+sky130_fd_pr__pfet_g5v0d16v0__vth0_diff_1+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d16v0__mm_mult*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope+0.0065)/sqrt(l*w*mult))'
+ k1 = 6.831000e-1
+ k2 = '-1.303200e-003+sky130_fd_pr__pfet_g5v0d16v0__k2_diff_1'
+ k3 = .000000e+0
+ k3b = .000000e+0
+ w0 = .000000e+0
+ dvt0 = .000000e+0
+ dvt1 = 5.300000e-1
+ dvt2 = -3.200000e-2
+ dvt0w = .000000e+0
+ dvt1w = 5.300000e+6
+ dvt2w = -3.200000e-2
+ dsub = '3.416000e-001+sky130_fd_pr__pfet_g5v0d16v0__dsub_diff_1'
+ minv = .000000e+0
+ voffl = .000000e+0
+ dvtp0 = .000000e+0
+ dvtp1 = .000000e+0
+ lpe0 = '1.400000e-007+sky130_fd_pr__pfet_g5v0d16v0__lpe0_diff_1'
+ lpeb = -6.500000e-8
+ vbm = -3.000000e+0
+ phin = .000000e+0
+ cdsc = 2.520000e-4
+ cdscb = .000000e+0
+ cdscd = .000000e+0
+ cit = .000000e+0
*(mismatch parameter sky130_fd_pr__pfet_g5v0d16v0__voff_slope_spectre)
+ voff = '-1.372000e-001+sky130_fd_pr__pfet_g5v0d16v0__voff_diff_1+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d16v0__mm_mult*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope+0.02)/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d16v0__nfactor_slope_spectre)
+ nfactor = '7.100000e-001+sky130_fd_pr__pfet_g5v0d16v0__nfactor_diff_1+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d16v0__mm_mult*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope+0.6)/sqrt(l*w*mult))'
+ eta0 = '8.729800e-002+sky130_fd_pr__pfet_g5v0d16v0__eta0_diff_1'
+ etab = -5.000000e-2
+ u0 = '2.707600e-002+sky130_fd_pr__pfet_g5v0d16v0__u0_diff_1'
+ ua = '2.585600e-009+sky130_fd_pr__pfet_g5v0d16v0__ua_diff_1'
+ ub = '4.595800e-019+sky130_fd_pr__pfet_g5v0d16v0__ub_diff_1'
+ uc = -1.220000e-10
+ eu = 1.670000e+0
+ vsat = '7.660800e+004+sky130_fd_pr__pfet_g5v0d16v0__vsat_diff_1'
+ a0 = '3.820000e-001+sky130_fd_pr__pfet_g5v0d16v0__a0_diff_1'
+ ags = '1.291200e-001+sky130_fd_pr__pfet_g5v0d16v0__ags_diff_1'
+ a1 = .000000e+0
+ a2 = 7.200000e-1
+ b0 = '4.000000e-012+sky130_fd_pr__pfet_g5v0d16v0__b0_diff_1'
+ b1 = '0.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__b1_diff_1'
+ keta = '-3.321800e-002+sky130_fd_pr__pfet_g5v0d16v0__keta_diff_1'
+ dwg = .000000e+0
+ dwb = .000000e+0
+ pclm = '1.000000e-001+sky130_fd_pr__pfet_g5v0d16v0__pclm_diff_1'
+ pdiblc1 = 3.900000e-1
+ pdiblc2 = 8.600000e-3
+ pdiblcb = -5.400000e-5
+ drout = 5.600000e-1
+ pvag = 5.040000e-1
+ delta = 8.900000e-3
+ pscbe1 = 5.088000e+8
+ pscbe2 = 6.945200e-9
+ fprout = .000000e+0
+ pdits = '0.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__pdits_diff_1'
+ pditsd = '0.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__pditsd_diff_1'
+ pditsl = .000000e+0
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = '3.310200e+002+sky130_fd_pr__pfet_g5v0d16v0__rdsw_diff_1'
+ rsw = 1.000000e+2
+ rdw = '1.000000e+001+sky130_fd_pr__pfet_g5v0d16v0__rdw_diff_1'
+ rdswmin = .000000e+0
+ rdwmin = .000000e+0
+ rswmin = .000000e+0
+ prwg = .000000e+0
+ prwb = -4.000000e-4
+ wr = 1.000000e+0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.000000e-7
+ alpha1 = 1.001000e+0
+ beta0 = 1.000000e+2
* Gidl Induced Drain Leakage Model Parameters
+ agidl = '1.650000e-010+sky130_fd_pr__pfet_g5v0d16v0__agidl_diff_1'
+ bgidl = '5.999300e+009+sky130_fd_pr__pfet_g5v0d16v0__bgidl_diff_1'
+ cgidl = '1.394000e+000+sky130_fd_pr__pfet_g5v0d16v0__cgidl_diff_1'
+ egidl = 4.920000e-2
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 1.160000e-8
+ aigbacc = '4.300000e-001+sky130_fd_pr__pfet_g5v0d16v0__aigbacc_diff_1'
+ bigbacc = 5.400000e-2
+ cigbacc = 7.500000e-2
+ nigbacc = '1.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__nigbacc_diff_1'
+ aigbinv = '3.500000e-001+sky130_fd_pr__pfet_g5v0d16v0__aigbinv_diff_1'
+ bigbinv = 3.000000e-2
+ cigbinv = 6.000000e-3
+ eigbinv = 1.100000e+0
+ nigbinv = '3.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__nigbinv_diff_1'
+ aigc = '4.300000e-001+sky130_fd_pr__pfet_g5v0d16v0__aigc_diff'
+ bigc = 5.400000e-2
+ cigc = 7.500000e-2
+ aigsd = '4.300000e-001+sky130_fd_pr__pfet_g5v0d16v0__aigsd_diff_1'
+ bigsd = '5.400000e-002+sky130_fd_pr__pfet_g5v0d16v0__bigsd_diff_1'
+ cigsd = 7.500000e-2
+ nigc = 1.000000e+0
+ poxedge = 1.000000e+0
+ pigcd = 1.000000e+0
+ ntox = 1.000000e+0
* Charge AND Capacitance Model Parameters
+ dlc = '-9.682600e-008+sky130_fd_pr__pfet_g5v0d16v0__dlc_diff+sky130_fd_pr__pfet_g5v0d16v0__dlc_rotweak'
+ dwc = '0.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__dwc_diff'
+ xpart = .000000e+0
+ cgso = '1.977100e-010*sky130_fd_pr__pfet_g5v0d16v0__soverlap_mult'
+ cgdo = '1.977100e-010*sky130_fd_pr__pfet_g5v0d16v0__doverlap_mult'
+ cgbo = .000000e+0
+ cgdl = '1.117200e-012*sky130_fd_pr__pfet_g5v0d16v0__doverlap_mult'
+ cgsl = '1.152000e-012*sky130_fd_pr__pfet_g5v0d16v0__soverlap_mult'
+ clc = 6.324000e-9
+ cle = 8.910000e-1
+ cf = '0.000000e+000+sky130_fd_pr__pfet_g5v0d16v0__cf_diff'
+ ckappas = 6.000000e-1
+ ckappad = 6.000000e-1
+ vfbcv = -1.000000e+0
+ acde = 9.129800e-1
+ moin = 1.556200e+1
+ noff = 1.045000e+0
+ voffcv = -1.815100e-1
* High-Speed/RF Model Parameters
* Flicker AND Thermal Noise Model Parameters
+ ef = 1.000000e+0
+ noia = 6.250000e+41
+ noib = 3.125000e+26
+ noic = 8.750000e+9
+ em = 4.100000e+7
* Layout-Dependent Parasitics Model Parameters
+ xl = .000000e+0
+ xw = .000000e+0
+ dmcg = .000000e+0
+ dmdg = .000000e+0
+ dmcgt = .000000e+0
+ xgw = .000000e+0
+ xgl = .000000e+0
+ ngcon = 1.000000e+0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.148300e-5
+ jsws = 4.020000e-12
+ jtssws = '4.020000e-012+sky130_fd_pr__pfet_g5v0d16v0__jtssws_diff_1'
+ ijthsfwd = 1.000000e-1
+ ijthsrev = 1.000000e-1
+ bvs = 1.269000e+1
+ xjbvs = 1.000000e+0
+ pbs = 6.587000e-1
+ cjs = '7.754700e-004*sky130_fd_pr__pfet_g5v0d16v0__ajunction_mult'
+ mjs = 3.395600e-1
+ pbsws = 1.000000e+0
+ cjsws = '9.871700e-011*sky130_fd_pr__pfet_g5v0d16v0__pjunction_mult'
+ mjsws = 2.467600e-1
+ pbswgs = 3.000000e+0
+ cjswgs = '1.460000e-010*sky130_fd_pr__pfet_g5v0d16v0__pjunction_mult'
+ mjswgs = 8.100000e-1
* Temperature Dependence Parameters
+ tnom = 3.000000e+1
+ kt1 = '-4.930800e-001+sky130_fd_pr__pfet_g5v0d16v0__kt1_diff_1'
+ kt1l = 1.000000e-11
+ kt2 = 5.633800e-4
+ ute = -1.646200e+0
+ ua1 = 1.218100e-9
+ ub1 = -1.241200e-18
+ uc1 = 8.272000e-12
+ prt = .000000e+0
+ at = -6.400000e+4
+ tvoff = '1.500000e-002+sky130_fd_pr__pfet_g5v0d16v0__tvoff_diff_1'
+ njs = 1.363200e+0
+ njd = 1.079100e+0
+ tpb = 1.671000e-3
+ tcj = 9.600000e-4
+ tpbsw = .000000e+0
+ tcjsw = 3.000000e-5
+ tpbswg = .000000e+0
+ tcjswg = .000000e+0
+ xtis = 1.000000e+1
+ xtid = 3.000000e+0
* DW AND DL Parameters
+ ll = .000000e+0
+ wl = .000000e+0
+ lln = 1.000000e+0
+ wln = 1.000000e+0
+ lw = .000000e+0
+ ww = .000000e+0
+ lwn = 1.000000e+0
+ wwn = 1.000000e+0
+ lwl = .000000e+0
+ wwl = .000000e+0
+ llc = .000000e+0
+ wlc = .000000e+0
+ lwc = .000000e+0
+ wwc = .000000e+0
+ lwlc = .000000e+0
+ wwlc = .000000e+0
* Stress Parameters
+ saref = .28e-6
+ sbref = 1.19e-6
+ kvth0 = '0.0+sky130_fd_pr__pfet_g5v0d16v0__kvth0_diff'
+ lkvth0 = '0.0+sky130_fd_pr__pfet_g5v0d16v0__lkvth0_diff'
+ wkvth0 = '0.0+sky130_fd_pr__pfet_g5v0d16v0__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 1.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0.0+sky130_fd_pr__pfet_g5v0d16v0__ku0_diff'
+ lku0 = '0.0+sky130_fd_pr__pfet_g5v0d16v0__lku0_diff'
+ wku0 = '0.0+sky130_fd_pr__pfet_g5v0d16v0__wku0_diff'
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 1.0
+ wlodku0 = 1.0
+ kvsat = '0.0+sky130_fd_pr__pfet_g5v0d16v0__kvsat_diff'
+ steta0 = 0.0
.ends sky130_fd_pr__pfet_g5v0d16v0__base
* Well Proximity Effect Parameters
