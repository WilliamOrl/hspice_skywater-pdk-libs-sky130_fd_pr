* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param GAU = AGAUSS(0,1.0,1)
* statistics '
* 	mismatch '
*     	'
*         process '
* 		vary sky130_fd_pr__res_xhigh_po__var_mult dist=gauss std=0.025
* 		vary sky130_fd_pr__res_high_po__var       dist=gauss std=0.025
*         '
* '
.subckt  sky130_fd_pr__res_xhigh_po__base r1 r2 b
+ 
+ w=1 l=1 mult=1
+ 
.param  rsheet = 2000.0
+ vc1_body = -1.00e-3
+ vc2_body = -1.00e-4
+ vc1_raw_end = -2.02e-2
+ vc2_raw_end = 1.55e-1
+ vc3_raw_end = 4.61e-2
+ body_pelgrom = 0.0347
+ r0_var = '17.23/w+2.318'
+ r1_var = '11.76/w'
+ rcon = '-46.62/(w*w)+331.73/w+20.576'
+ rend_mm = '0.0472/sqrt(w)'
+ tc1_voltco = -7.1e-3
+ rend_var = 'sky130_fd_pr__res_high_po__var_mult*sqrt(2)*r0_var'
+ rtot_var = 'sky130_fd_pr__res_high_po__var_mult*sqrt(2*pow(r0_var,2)+pow((r1_var*l),2))'
*(mismatch parameter sky130_fd_pr__res_high_po__slope_spectre)
+ res_match = '(body_pelgrom/sqrt(w*l*mult))*MC_MM_SWITCH*GAU'
+ rbody_var = 'rtot_var-rend_var'
*(mismatch parameter sky130_fd_pr__res_high_po__con_slope_spectre)
+ rend = '(rcon+rend_var)*(1+rend_mm/sqrt(mult)*MC_MM_SWITCH*GAU)'
+ vc1_end = 'vc1_raw_end/pwr(l,0.5)*(1+tc1_voltco*(temper-30))'
+ vc2_end = 'vc2_raw_end/pwr(l,0.5)*(1+tc1_voltco*(temper-30))'
+ vc3_end = 'vc3_raw_end/pwr(l,0.5)*(1+tc1_voltco*(temper-30))'
+ rbody = '(l*rsheet+rbody_var)*(1+res_match)/w'
rbody ra r2 r = 'rbody*(1+abs(v(r1,r2))*vc1_body+abs(v(r1,r2))*abs(v(r1,r2))/(l*l)*vc2_body)'
+ tc1 = -1.47e-3
+ tc2 = 2.7e-6
*+tnom = 30.0
rend r1 ra  r = 'rend*(1+vc1_raw_end*(1-exp(-abs(v(r2,r1))))+
+ vc2_raw_end*(1 - exp(-abs(v(r2,r1)))) * (1 - exp(-abs(v(r2,r1)))) +
+ vc3_raw_end*(1 - exp(-abs(v(r2,r1)))) * (1 - exp(-abs(v(r2,r1)))) * (1 - exp(-abs(v(r2,r1))))       ) '
c1 r2 b  c = '((l+2*2.08)*w*crpf_precision*1e-12+2*(l+2*2.08+w)*crpfsw_precision_1_1*1e-6)/2'
c2 r1 b  c = '((l+2*2.08)*w*crpf_precision*1e-12+2*(l+2*2.08+w)*crpfsw_precision_1_1*1e-6)/2'
.ends sky130_fd_pr__res_xhigh_po__base
