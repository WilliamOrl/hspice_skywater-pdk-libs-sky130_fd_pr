* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.subckt  sky130_fd_pr__esd_nfet_01v8 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__esd_nfet_01v8 d g s b sky130_fd_pr__esd_nfet_01v8__model l = 'l' w = 'w' nf = 'nf' ad = 'ad' as = 'as' pd = 'pd' ps = 'ps' nrd = 'nrd' nrs = 'nrs' sa = 'sa' sb = 'sb' sd = 'sd'
.model sky130_fd_pr__esd_nfet_01v8__model.0 nmos
* DC IV MOS Parameters
+ lmin = 1.6e-07 lmax = 1.7e-07 wmin = 2.0345e-05 wmax = 2.0355e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.1482e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '1.2561e-008+sky130_fd_pr__esd_nfet_01v8__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '1.1879846e-008+sky130_fd_pr__esd_nfet_01v8__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 200000.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.1482e-009*sky130_fd_pr__esd_nfet_01v8__toxe_mult'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__esd_nfet_01v8__rshn_mult'
* Threshold Voltage Parameters
+ vth0 = '0.565+sky130_fd_pr__esd_nfet_01v8__vth0_diff_0'
+ k1 = 0.50824
+ k2 = '-0.036074+sky130_fd_pr__esd_nfet_01v8__k2_diff_0'
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 8.8387e-8
+ lpeb = -7.1972e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '163960+sky130_fd_pr__esd_nfet_01v8__vsat_diff_0'
+ ua = '-1.244e-009+sky130_fd_pr__esd_nfet_01v8__ua_diff_0'
+ ub = '1.6282e-018+sky130_fd_pr__esd_nfet_01v8__ub_diff_0'
+ uc = 1.9958e-11
+ rdsw = '174.5+sky130_fd_pr__esd_nfet_01v8__rdsw_diff_0'
+ prwb = -0.17995
+ prwg = 0.011
+ wr = 1.0
+ u0 = '0.028432+sky130_fd_pr__esd_nfet_01v8__u0_diff_0'
+ a0 = '1.5+sky130_fd_pr__esd_nfet_01v8__a0_diff_0'
+ keta = '0.0873+sky130_fd_pr__esd_nfet_01v8__keta_diff_0'
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = '0.4092+sky130_fd_pr__esd_nfet_01v8__ags_diff_0'
+ b0 = '0+sky130_fd_pr__esd_nfet_01v8__b0_diff_0'
+ b1 = '0+sky130_fd_pr__esd_nfet_01v8__b1_diff_0'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1848+sky130_fd_pr__esd_nfet_01v8__voff_diff_0'
+ nfactor = '2+sky130_fd_pr__esd_nfet_01v8__nfactor_diff_0'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = '0+sky130_fd_pr__esd_nfet_01v8__tvoff_diff_0'
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = '0+sky130_fd_pr__esd_nfet_01v8__eta0_diff_0'
+ etab = 0.001
+ dsub = 0.1
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = '0.17122+sky130_fd_pr__esd_nfet_01v8__pclm_diff_0'
+ pdiblc1 = 0.10049528
+ pdiblc2 = 0.020103
+ pdiblcb = -1.0
+ drout = 0.48621
+ pscbe1 = 3.6928e+8
+ pscbe2 = 2.2e-6
+ pvag = 0.0
+ delta = 0.01184
+ alpha0 = 1.414e-6
+ alpha1 = 1.4744
+ beta0 = 17.6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '3.041136e-013+sky130_fd_pr__esd_nfet_01v8__pdits_diff_0'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__esd_nfet_01v8__pditsd_diff_0'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.1482e-9
* Temperature Effects Parameters
+ kt1 = '-0.29744+sky130_fd_pr__esd_nfet_01v8__kt1_diff_0'
+ kt2 = -0.019143
+ at = 79266.0
+ ute = -1.6806
+ ua1 = 5.504e-10
+ ub1 = 2.7351e-19
+ uc1 = 1.6706e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = '3.2e-010*sky130_fd_pr__esd_nfet_01v8__overlap_mult'
+ cgso = '3.2e-010*sky130_fd_pr__esd_nfet_01v8__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__esd_nfet_01v8__overlap_mult'
+ cgdl = '0*sky130_fd_pr__esd_nfet_01v8__overlap_mult'
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = '1.8739e-008+sky130_fd_pr__esd_nfet_01v8__dlc_diff+sky130_fd_pr__esd_nfet_01v8__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__esd_nfet_01v8__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.621
+ voffcv = -0.1372
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.0013459*sky130_fd_pr__esd_nfet_01v8__ajunction_mult'
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = '3.6001e-011*sky130_fd_pr__esd_nfet_01v8__pjunction_mult'
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = '2.3347e-010*sky130_fd_pr__esd_nfet_01v8__pjunction_mult'
+ mjswgs = 0.8000
+ pbswgs = 0.95578
.model sky130_fd_pr__esd_nfet_01v8__model.1 nmos
* DC IV MOS Parameters
+ lmin = 1.6e-07 lmax = 1.7e-07 wmin = 4.0305e-05 wmax = 4.0315e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.1482e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '1.2561e-008+sky130_fd_pr__esd_nfet_01v8__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '1.1879846e-008+sky130_fd_pr__esd_nfet_01v8__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 200000.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.1482e-009*sky130_fd_pr__esd_nfet_01v8__toxe_mult'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__esd_nfet_01v8__rshn_mult'
* Threshold Voltage Parameters
+ vth0 = '0.574+sky130_fd_pr__esd_nfet_01v8__vth0_diff_1'
+ k1 = 0.47947
+ k2 = '-0.0071285+sky130_fd_pr__esd_nfet_01v8__k2_diff_1'
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 8.8387e-8
+ lpeb = -7.1972e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '162130+sky130_fd_pr__esd_nfet_01v8__vsat_diff_1'
+ ua = '-1.3196e-009+sky130_fd_pr__esd_nfet_01v8__ua_diff_1'
+ ub = '1.5781e-018+sky130_fd_pr__esd_nfet_01v8__ub_diff_1'
+ uc = 1.9293e-11
+ rdsw = '174.5+sky130_fd_pr__esd_nfet_01v8__rdsw_diff_1'
+ prwb = -0.17995
+ prwg = 0.011
+ wr = 1.0
+ u0 = '0.028739+sky130_fd_pr__esd_nfet_01v8__u0_diff_1'
+ a0 = '1.5+sky130_fd_pr__esd_nfet_01v8__a0_diff_1'
+ keta = '0.072913+sky130_fd_pr__esd_nfet_01v8__keta_diff_1'
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = '0.4092+sky130_fd_pr__esd_nfet_01v8__ags_diff_1'
+ b0 = '0+sky130_fd_pr__esd_nfet_01v8__b0_diff_1'
+ b1 = '0+sky130_fd_pr__esd_nfet_01v8__b1_diff_1'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1936+sky130_fd_pr__esd_nfet_01v8__voff_diff_1'
+ nfactor = '2+sky130_fd_pr__esd_nfet_01v8__nfactor_diff_1'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = '0+sky130_fd_pr__esd_nfet_01v8__tvoff_diff_1'
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = '0+sky130_fd_pr__esd_nfet_01v8__eta0_diff_1'
+ etab = 0.001
+ dsub = 0.1
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = '0.15544+sky130_fd_pr__esd_nfet_01v8__pclm_diff_1'
+ pdiblc1 = 0.10049528
+ pdiblc2 = 0.030979
+ pdiblcb = -1.0
+ drout = 0.57882
+ pscbe1 = 3.6928e+8
+ pscbe2 = 2.2e-6
+ pvag = 0.0
+ delta = 0.01376
+ alpha0 = 1.414e-6
+ alpha1 = 1.4744
+ beta0 = 17.6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '3.041136e-013+sky130_fd_pr__esd_nfet_01v8__pdits_diff_1'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__esd_nfet_01v8__pditsd_diff_1'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.1482e-9
* Temperature Effects Parameters
+ kt1 = '-0.29351+sky130_fd_pr__esd_nfet_01v8__kt1_diff_1'
+ kt2 = -0.019143
+ at = 71264.0
+ ute = -1.6806
+ ua1 = 5.7242e-10
+ ub1 = 9.1861e-19
+ uc1 = 1.6038e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = '3.2e-010*sky130_fd_pr__esd_nfet_01v8__overlap_mult'
+ cgso = '3.2e-010*sky130_fd_pr__esd_nfet_01v8__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__esd_nfet_01v8__overlap_mult'
+ cgdl = '0*sky130_fd_pr__esd_nfet_01v8__overlap_mult'
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = '1.8739e-008+sky130_fd_pr__esd_nfet_01v8__dlc_diff+sky130_fd_pr__esd_nfet_01v8__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__esd_nfet_01v8__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.621
+ voffcv = -0.1372
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.0013459*sky130_fd_pr__esd_nfet_01v8__ajunction_mult'
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = '3.6001e-011*sky130_fd_pr__esd_nfet_01v8__pjunction_mult'
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = '2.3347e-010*sky130_fd_pr__esd_nfet_01v8__pjunction_mult'
+ mjswgs = 0.8000
+ pbswgs = 0.95578
.model sky130_fd_pr__esd_nfet_01v8__model.2 nmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 5.395e-06 wmax = 5.405e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.1482e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '1.2561e-008+sky130_fd_pr__esd_nfet_01v8__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '1.1879846e-008+sky130_fd_pr__esd_nfet_01v8__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 200000.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.1482e-009*sky130_fd_pr__esd_nfet_01v8__toxe_mult'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__esd_nfet_01v8__rshn_mult'
* Threshold Voltage Parameters
+ vth0 = '0.59966+sky130_fd_pr__esd_nfet_01v8__vth0_diff_2'
+ k1 = 0.47947
+ k2 = '-0.008+sky130_fd_pr__esd_nfet_01v8__k2_diff_2'
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 8.8387e-8
+ lpeb = -7.1972e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '140380+sky130_fd_pr__esd_nfet_01v8__vsat_diff_2'
+ ua = '-1.1107e-009+sky130_fd_pr__esd_nfet_01v8__ua_diff_2'
+ ub = '1.6158e-018+sky130_fd_pr__esd_nfet_01v8__ub_diff_2'
+ uc = 3.08e-11
+ rdsw = '174.5+sky130_fd_pr__esd_nfet_01v8__rdsw_diff_2'
+ prwb = -0.17995
+ prwg = 0.011
+ wr = 1.0
+ u0 = '0.029546+sky130_fd_pr__esd_nfet_01v8__u0_diff_2'
+ a0 = '1.5+sky130_fd_pr__esd_nfet_01v8__a0_diff_2'
+ keta = '0.0873+sky130_fd_pr__esd_nfet_01v8__keta_diff_2'
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = '0.4092+sky130_fd_pr__esd_nfet_01v8__ags_diff_2'
+ b0 = '0+sky130_fd_pr__esd_nfet_01v8__b0_diff_2'
+ b1 = '0+sky130_fd_pr__esd_nfet_01v8__b1_diff_2'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1936+sky130_fd_pr__esd_nfet_01v8__voff_diff_2'
+ nfactor = '2+sky130_fd_pr__esd_nfet_01v8__nfactor_diff_2'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = '0+sky130_fd_pr__esd_nfet_01v8__tvoff_diff_2'
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = '0.00078661337+sky130_fd_pr__esd_nfet_01v8__eta0_diff_2'
+ etab = -0.0029133829
+ dsub = 0.1
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = '0.33234+sky130_fd_pr__esd_nfet_01v8__pclm_diff_2'
+ pdiblc1 = 0.10049528
+ pdiblc2 = 0.015545
+ pdiblcb = -1.0
+ drout = 0.87701
+ pscbe1 = 3.6928e+8
+ pscbe2 = 2.0e-6
+ pvag = 0.0
+ delta = 0.008
+ alpha0 = 1.414e-6
+ alpha1 = 1.4744
+ beta0 = 17.6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '3.041136e-013+sky130_fd_pr__esd_nfet_01v8__pdits_diff_2'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__esd_nfet_01v8__pditsd_diff_2'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.1482e-9
* Temperature Effects Parameters
+ kt1 = '-0.33011+sky130_fd_pr__esd_nfet_01v8__kt1_diff_2'
+ kt2 = -0.019143
+ at = 77739.0
+ ute = -1.6806
+ ua1 = 5.504e-10
+ ub1 = 4.8841e-19
+ uc1 = 1.6706e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = '3.2e-010*sky130_fd_pr__esd_nfet_01v8__overlap_mult'
+ cgso = '3.2e-010*sky130_fd_pr__esd_nfet_01v8__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__esd_nfet_01v8__overlap_mult'
+ cgdl = '0*sky130_fd_pr__esd_nfet_01v8__overlap_mult'
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = '1.8739e-008+sky130_fd_pr__esd_nfet_01v8__dlc_diff+sky130_fd_pr__esd_nfet_01v8__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__esd_nfet_01v8__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.621
+ voffcv = -0.1372
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.0013459*sky130_fd_pr__esd_nfet_01v8__ajunction_mult'
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = '3.6001e-011*sky130_fd_pr__esd_nfet_01v8__pjunction_mult'
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = '2.3347e-010*sky130_fd_pr__esd_nfet_01v8__pjunction_mult'
+ mjswgs = 0.8000
+ pbswgs = 0.95578
.ends sky130_fd_pr__esd_nfet_01v8
