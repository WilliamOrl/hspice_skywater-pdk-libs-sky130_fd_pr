* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* ./parameters_cap_nom.spice created from ./parameters.spice
*
.param GAU = AGAUSS(0,0.0475,1)
.param GAU2 = AGAUSS(0,0.1,1)
.param GAU3 = AGAUSS(0,2.4e-08,1)

.param sw_fox_cap = '1.0+corner_factor*0.0' + process_mc_factor*MC_PR_SWITCH*GAU
.param sw_fox_poly_cap = '1.0+corner_factor*0.0' + process_mc_factor*MC_PR_SWITCH*GAU
.param sw_li_cap = '1.0+corner_factor*0.0' + process_mc_factor*MC_PR_SWITCH*EXP(GAU2)
.param sw_cap_mim_ca = '2e-15+corner_factor*0.0' + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.027000000000000003,1)
.param sw_cap_mim_dw = '1.5e-07+corner_factor*0.0' + process_mc_factor*MC_PR_SWITCH*GAU3
