* SKY130 Spice File.
* Slow    Varactor Parameters
.param
+ cnwvc_tox='41.6503*1.024*1.06'
+ cnwvc_cdepmult=0.9
+ cnwvc_cintmult=0.95
+ cnwvc_vt1='0.3333+0.112'
+ cnwvc_vt2='0.2380952+0.112'
+ cnwvc_vtr='0.16+0.112'
+ cnwvc_dwc=-0.02
+ cnwvc_dlc=-0.01
+ cnwvc_dld=-0.0008
+ cnwvc2_tox='41.7642*1.017*1.06'
+ cnwvc2_cdepmult=0.95
+ cnwvc2_cintmult=0.95
+ cnwvc2_vt1='0.2+0.074'
+ cnwvc2_vt2='0.33+0.074'
+ cnwvc2_vtr='0.14+0.074'
+ cnwvc2_dwc=-0.02
+ cnwvc2_dlc=-0.01
+ cnwvc2_dld=-0.0006
* sky130_fd_pr__model__parasitic__diode_ps2nw Parameters
.param
+ sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult = 1.1178e+00    
+ sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult = 1.0401e+00    
* sky130_fd_pr__model__parasitic__diode_ps2dn Parameters
+ sky130_fd_pr__model__parasitic__diode_ps2dn__ajunction_mult = 1.174      
+ sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult = 1.234       
* sky130_fd_pr__model__parasitic__diode_pw2dn Parameters
+ sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult = 1.189    
+ sky130_fd_pr__model__parasitic__diode_pw2dn__pjunction_mult = 1.008    
* sky130_fd_pr__diode_pw2nd_05v5  Parameters
+ sky130_fd_pr__nfet_01v8__ajunction_mult = 1.1505e+0
+ sky130_fd_pr__nfet_01v8__pjunction_mult = 1.1793e+0
* sky130_fd_pr__diode_pd2nw_05v5_hvt  Parameters
+ sky130_fd_pr__pfet_01v8_hvt__ajunction_mult = 1.0491e+0
+ sky130_fd_pr__pfet_01v8_hvt__pjunction_mult = 1.0970e+0
+ dkispp=7.0967e-01 dkbfpp=4.9061e-01 dknfpp=1.000
+ dkispp5x=7.8658e-01 dkbfpp5x=4.6158e-01 dknfpp5x=1.0009e+00 dkisepp5x=0.745
+ cvpp2_nhvnative10x4_cor=0.862
+ cvpp2_nhvnative10x4_sub=8.68e-16
+ cvpp2_phv5x4_cor=0.862
+ cvpp2_phv5x4_sub=8.68e-16
