* Copyright 2022 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SKY130 Spice File.
* Critical Model Parameters:
.param GAU = AGAUSS(0,1.0,1)
.param GAU2 = AGAUSS(0,1.5,1)
.param GAU3 = AGAUSS(0,2.8,1)
.param GAU4 = AGAUSS(0,0.8,1)
.param GAU5 = AGAUSS(0,0.6,1)
.param GAU6 = AGAUSS(0,1.8,1)
.param GAU7 = AGAUSS(0,2.0,1)
.param GAU8 = AGAUSS(0,1.1,1)
.param GAU9 = AGAUSS(0,0.5,1)
.param GAU10 = AGAUSS(0,0.3,1)
.param GAU11 = AGAUSS(0,1.3,1)

.param cnwvc = 0.0 + MC_PR_SWITCH*GAU
.param diff_cd = 0.0 + MC_PR_SWITCH*GAU2
.param hvn_bodyeffect = 0.0 + MC_PR_SWITCH*GAU3
.param hvn_diode = 0.0 + MC_PR_SWITCH*GAU
.param hvn_mobility = 0.0 + MC_PR_SWITCH*GAU4
.param hvn_saturation = 0.0 + MC_PR_SWITCH*GAU5
.param hvn_subvt = 0.0 + MC_PR_SWITCH*GAU
.param hvn_threshold = 0.0 + MC_PR_SWITCH*GAU2
.param hvp_bodyeffect = 0.0 + MC_PR_SWITCH*GAU3
.param hvp_diode = 0.0 + MC_PR_SWITCH*GAU
.param hvp_mobility = 0.0 + MC_PR_SWITCH*GAU6
.param hvp_saturation = 0.0 + MC_PR_SWITCH*GAU6
.param hvp_subvt = 0.0 + MC_PR_SWITCH*GAU
.param hvp_threshold = 0.0 + MC_PR_SWITCH*GAU2
.param hvtox = 0.0 + MC_PR_SWITCH*GAU
.param ic_cap = 0.0 + MC_PR_SWITCH*GAU
.param ic_res = 0.0 + MC_PR_SWITCH*GAU
.param ic_res_ndiff = 0.0 + MC_PR_SWITCH*GAU
.param ic_res_pdiff = 0.0 + MC_PR_SWITCH*GAU
.param ic_res_poly = 0.0 + MC_PR_SWITCH*GAU
.param ic_res_pwell = 0.0 + MC_PR_SWITCH*GAU
.param lvhp_bodyeffect = 0.0 + MC_PR_SWITCH*GAU6
.param lvhp_mobility = 0.0 + MC_PR_SWITCH*GAU7
.param lvhp_saturation = 0.0 + MC_PR_SWITCH*GAU8
.param lvhp_threshold = 0.0 + MC_PR_SWITCH*GAU4
.param lvln_bodyeffect = 0.0 + MC_PR_SWITCH*GAU7
.param lvln_mobility = 0.0 + MC_PR_SWITCH*GAU5
.param lvln_saturation = 0.0 + MC_PR_SWITCH*GAU5
.param lvln_threshold = 0.0 + MC_PR_SWITCH*GAU5
.param lvlp_bodyeffect = 0.0 + MC_PR_SWITCH*GAU9
.param lvlp_mobility = 0.0 + MC_PR_SWITCH*GAU10
.param lvlp_saturation = 0.0 + MC_PR_SWITCH*GAU10
.param lvlp_threshold = 0.0 + MC_PR_SWITCH*GAU11
.param lvn_bodyeffect = 0.0 + MC_PR_SWITCH*GAU7
.param lvn_diode = 0.0 + MC_PR_SWITCH*GAU
.param lvn_mobility = 0.0 + MC_PR_SWITCH*GAU5
.param lvn_saturation = 0.0 + MC_PR_SWITCH*GAU5
.param lvn_subvt = 0.0 + MC_PR_SWITCH*GAU
.param lvn_threshold = 0.0 + MC_PR_SWITCH*GAU4
.param lvp_bodyeffect = 0.0 + MC_PR_SWITCH*GAU
.param lvp_diode = 0.0 + MC_PR_SWITCH*GAU
.param lvp_mobility = 0.0 + MC_PR_SWITCH*GAU7
.param lvp_saturation = 0.0 + MC_PR_SWITCH*GAU8
.param lvp_subvt = 0.0 + MC_PR_SWITCH*GAU
.param lvp_threshold = 0.0 + MC_PR_SWITCH*GAU
.param lvtox = 0.0 + MC_PR_SWITCH*GAU8
.param mim = 0.0 + MC_PR_SWITCH*GAU
.param hvntvn_threshold = 0.0 + MC_PR_SWITCH*GAU
.param nfet_20v0_nvt = 0.0 + MC_PR_SWITCH*GAU
.param nfet_20v0_nvt_iso = 0.0 + MC_PR_SWITCH*GAU
.param nfet_20v0 = 0.0 + MC_PR_SWITCH*GAU
.param nfet_20v0_iso = 0.0 + MC_PR_SWITCH*GAU
.param n20zvtvh1defet = 0.0 + MC_PR_SWITCH*GAU
.param nfet_20v0_zvt = 0.0 + MC_PR_SWITCH*GAU
.param ndiff_cd = 0.0 + MC_PR_SWITCH*GAU2
.param pfet_20v0 = 0.0 + MC_PR_SWITCH*GAU
.param pdiff_cd = 0.0 + MC_PR_SWITCH*GAU2
.param nfet_01v8_lvt = 0.0 + MC_PR_SWITCH*GAU
.param special_nfet_pass_lvt = 0.0 + MC_PR_SWITCH*GAU
.param sky130_fd_pr__npn_05v5_all = 0.0 + MC_PR_SWITCH*GAU
.param nfet_g5v0d16v0 = 0.0 + MC_PR_SWITCH*GAU
.param pfet_01v8_mvt = 0.0 + MC_PR_SWITCH*GAU
.param pnp_05v5_W0p68L0p68 = 0.0 + MC_PR_SWITCH*GAU
.param poly_cd = 0.0 + MC_PR_SWITCH*GAU2
.param pfet_01v8 = 0.0 + MC_PR_SWITCH*GAU
.param pfet_g5v0d16v0 = 0.0 + MC_PR_SWITCH*GAU
.param well_diode = 0.0 + MC_PR_SWITCH*GAU
* statistics '
*  process '
*     vary cnwvc dist=gauss std=1.0
*     vary diff_cd dist=gauss std=1.5
*     vary hvn_bodyeffect dist=gauss std=2.8
*     vary hvn_diode dist=gauss std=1.0
*     vary hvn_mobility dist=gauss std=0.8
*     vary hvn_saturation dist=gauss std=0.6
*     vary hvn_subvt dist=gauss std=1.0
*     vary hvn_threshold dist=gauss std=1.5
*     vary hvp_bodyeffect dist=gauss std=2.8
*     vary hvp_diode dist=gauss std=1.0
*     vary hvp_mobility dist=gauss std=1.8
*     vary hvp_saturation dist=gauss std=1.8
*     vary hvp_subvt dist=gauss std=1.0
*     vary hvp_threshold dist=gauss std=1.5
*     vary hvtox dist=gauss std=1.0
*     vary ic_cap dist=gauss std=1.0
*     vary ic_res dist=gauss std=1.0
*     vary ic_res_ndiff dist=gauss std=1.0
*     vary ic_res_pdiff dist=gauss std=1.0
*     vary ic_res_poly dist=gauss std=1.0
*     vary ic_res_pwell dist=gauss std=1.0
*     vary lvhp_bodyeffect dist=gauss std=1.8
*     vary lvhp_mobility dist=gauss std=2.0
*     vary lvhp_saturation dist=gauss std=1.1
*     vary lvhp_threshold dist=gauss std=0.8
*     vary lvln_bodyeffect dist=gauss std=2.0
*     vary lvln_mobility dist=gauss std=0.6
*     vary lvln_saturation dist=gauss std=0.6
*     vary lvln_threshold dist=gauss std=0.6
*     vary lvlp_bodyeffect dist=gauss std=0.5
*     vary lvlp_mobility dist=gauss std=0.3
*     vary lvlp_saturation dist=gauss std=0.3
*     vary lvlp_threshold dist=gauss std=1.3
*     vary lvn_bodyeffect dist=gauss std=2.0
*     vary lvn_diode dist=gauss std=1.0
*     vary lvn_mobility dist=gauss std=0.6
*     vary lvn_saturation dist=gauss std=0.6
*     vary lvn_subvt dist=gauss std=1.0
*     vary lvn_threshold dist=gauss std=0.8
*     vary lvp_bodyeffect dist=gauss std=1.0
*     vary lvp_diode dist=gauss std=1.0
*     vary lvp_mobility dist=gauss std=2.0
*     vary lvp_saturation dist=gauss std=1.1
*     vary lvp_subvt dist=gauss std=1.0
*     vary lvp_threshold dist=gauss std=1.0
*     vary lvtox dist=gauss std=1.1
*     vary mim dist=gauss std=1.0
*     vary hvntvn_threshold dist=gauss std=1.0
*     vary nfet_20v0_nvt dist=gauss std=1.0
*     vary nfet_20v0_nvt_iso dist=gauss std=1.0
*     vary nfet_20v0 dist=gauss std=1.0
*     vary nfet_20v0_iso dist=gauss std=1.0
*     vary n20zvtvh1defet dist=gauss std=1.0
*     vary nfet_20v0_zvt dist=gauss std=1.0
*     vary ndiff_cd dist=gauss std=1.5
*     vary pfet_20v0 dist=gauss std=1.0
*     vary pdiff_cd dist=gauss std=1.5
*     vary nfet_01v8_lvt dist=gauss std=1.0
*     vary special_nfet_pass_lvt dist=gauss std=1.0
*     vary sky130_fd_pr__npn_05v5_all dist=gauss std=1.0
*     vary nfet_g5v0d16v0 dist=gauss std=1.0
*     vary pfet_01v8_mvt dist=gauss std=1.0
*     vary pnp_05v5_W0p68L0p68 dist=gauss std=1.0
*     vary poly_cd dist=gauss std=1.5
*     vary pfet_01v8 dist=gauss std=1.0
*     vary pfet_g5v0d16v0 dist=gauss std=1.0
*     vary well_diode dist=gauss std=1.0
*   '
*   mismatch '
*   '
* '
