* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param GAU = AGAUSS(0,1.0,1)
.param sky130_fd_pr__esd_nfet_05v0_nvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__esd_nfet_05v0_nvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__esd_nfet_05v0_nvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__esd_nfet_05v0_nvt__nfactor_slope_spectre = 0.0
* statistics '
*   process '
*   '
*   mismatch '
*     vary sky130_fd_pr__esd_nfet_05v0_nvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__esd_nfet_05v0_nvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__esd_nfet_05v0_nvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__esd_nfet_05v0_nvt__nfactor_slope_spectre dist=gauss std = 1.0
*   '
* '
.subckt  sky130_fd_pr__esd_nfet_05v0_nvt d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__esd_nfet_05v0_nvt d g s b sky130_fd_pr__esd_nfet_05v0_nvt__model l = 'l' w = 'w' nf = 'nf' ad = 'ad' as = 'as' pd = 'pd' ps = 'ps' nrd = 'nrd' nrs = 'nrs' sa = 'sa' sb = 'sb' sd = 'sd'
.model sky130_fd_pr__esd_nfet_05v0_nvt__model.0 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 9.995e-06 wmax = 1.0005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '6.93e-008+sky130_fd_pr__nfet_05v0_nvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '4.5e-008+sky130_fd_pr__nfet_05v0_nvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.6e-9
+ dwb = 1.92e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.8
+ rnoib = 0.38
+ tnoia = 7.6e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__esd_nfet_05v0_nvt__toxe_slope_spectre)
+ toxe = '1.16e-008*sky130_fd_pr__nfet_05v0_nvt__toxe_mult+MC_MM_SWITCH*GAU*(1.16e-008*sky130_fd_pr__nfet_05v0_nvt__toxe_mult*(sky130_fd_pr__nfet_05v0_nvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__nfet_05v0_nvt__rshn_mult'
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__esd_nfet_05v0_nvt__vth0_slope_spectre)
+ vth0 = '0.053+sky130_fd_pr__nfet_05v0_nvt__vth0_diff_0+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_05v0_nvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.364
+ k2 = '0.038817+sky130_fd_pr__nfet_05v0_nvt__k2_diff_0'
+ k3 = 1.4
+ dvt0 = 5.7
+ dvt1 = 0.21851
+ dvt2 = 0.04
+ dvt0w = 7.7
+ dvt1w = 1272000.0
+ dvt2w = -0.032
+ w0 = 0.0
+ k3b = -0.58
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = -1.2362266e-14
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '68940+sky130_fd_pr__nfet_05v0_nvt__vsat_diff_0'
+ ua = '8.4094e-010+sky130_fd_pr__nfet_05v0_nvt__ua_diff_0'
+ ub = '1.2863e-018+sky130_fd_pr__nfet_05v0_nvt__ub_diff_0'
+ uc = 3.2583e-11
+ rdsw = '430+sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_0'
+ prwb = 0.0
+ prwg = 1.0e-12
+ wr = 1.0
+ u0 = '0.050801+sky130_fd_pr__nfet_05v0_nvt__u0_diff_0'
+ a0 = '0.08+sky130_fd_pr__nfet_05v0_nvt__a0_diff_0'
+ keta = '-0.019904+sky130_fd_pr__nfet_05v0_nvt__keta_diff_0'
+ a1 = 0.0
+ a2 = 0.96293372
+ ags = '0.87995+sky130_fd_pr__nfet_05v0_nvt__ags_diff_0'
+ b0 = '3.3993e-007+sky130_fd_pr__nfet_05v0_nvt__b0_diff_0'
+ b1 = '0+sky130_fd_pr__nfet_05v0_nvt__b1_diff_0'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__esd_nfet_05v0_nvt__voff_slope_spectre)
+ voff = '0+sky130_fd_pr__nfet_05v0_nvt__voff_diff_0+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_05v0_nvt__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__esd_nfet_05v0_nvt__nfactor_slope_spectre)
+ nfactor = '0.63313+sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_0+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_05v0_nvt__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = '0+sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_0'
+ cit = 9.2584123e-8
+ cdsc = 0.0
+ cdscb = 1.4150948e-7
+ cdscd = 1.5e-5
+ eta0 = '9+sky130_fd_pr__nfet_05v0_nvt__eta0_diff_0'
+ etab = -0.00021692
+ dsub = 0.42
* BSIM4 - Sub-threshold parameters
+ voffl = 1.9445332e-8
+ minv = 0.0
* Rout Parameters
+ pclm = '0.11748+sky130_fd_pr__nfet_05v0_nvt__pclm_diff_0'
+ pdiblc1 = 8.833e-7
+ pdiblc2 = 0.0002
+ pdiblcb = 0.0
+ drout = 0.13139
+ pscbe1 = 2.4476e+8
+ pscbe2 = 3.84e-9
+ pvag = 4.5419436
+ delta = 0.007
+ alpha0 = 2.0236e-6
+ alpha1 = 0.093632
+ beta0 = 22.1
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0.02+sky130_fd_pr__nfet_05v0_nvt__pdits_diff_0'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_0'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = '-0.35858+sky130_fd_pr__nfet_05v0_nvt__kt1_diff_0'
+ kt2 = -0.016016
+ at = 11600.0
+ ute = -1.7861
+ ua1 = 4.4e-10
+ ub1 = -1.4256e-18
+ uc1 = -3.94e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.5764
+ jss = 0.00042966
+ jsws = 8.040000000000001e-10
+ xtis = 0.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019685
+ tpbsw = 0.001
+ tpbswg = 0.0
+ tcj = 0.00083
+ tcjsw = 0.0
+ tcjswg = 0.0
+ cgdo = '3.473e-010*sky130_fd_pr__nfet_05v0_nvt__overlap_mult'
+ cgso = '3.473e-010*sky130_fd_pr__nfet_05v0_nvt__overlap_mult'
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '5e-011*sky130_fd_pr__nfet_05v0_nvt__overlap_mult'
+ cgdl = '5e-011*sky130_fd_pr__nfet_05v0_nvt__overlap_mult'
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = '7.6493e-008+sky130_fd_pr__nfet_05v0_nvt__dlc_diff+sky130_fd_pr__nfet_05v0_nvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__nfet_05v0_nvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 1.16
+ moin = 15.0
+ noff = 4.0
+ voffcv = 0.216
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.0008602*sky130_fd_pr__nfet_05v0_nvt__ajunction_mult'
+ mjs = 0.28329
+ pbs = 0.66345
+ cjsws = '8.5152e-011*sky130_fd_pr__nfet_05v0_nvt__pjunction_mult'
+ mjsws = 0.057926
+ pbsws = 1.0
+ cjswgs = '3.58e-011*sky130_fd_pr__nfet_05v0_nvt__pjunction_mult'
+ mjswgs = 0.33
+ pbswgs = 0.2442
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__nfet_05v0_nvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__nfet_05v0_nvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__nfet_05v0_nvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__nfet_05v0_nvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__nfet_05v0_nvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__nfet_05v0_nvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__nfet_05v0_nvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__nfet_05v0_nvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__esd_nfet_05v0_nvt__model.1 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 9.995e-06 wmax = 1.0005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '6.93e-008+sky130_fd_pr__nfet_05v0_nvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '4.5e-008+sky130_fd_pr__nfet_05v0_nvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.6e-9
+ dwb = 1.92e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.8
+ rnoib = 0.38
+ tnoia = 7.6e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__esd_nfet_05v0_nvt__toxe_slope_spectre)
+ toxe = '1.16e-008*sky130_fd_pr__nfet_05v0_nvt__toxe_mult+MC_MM_SWITCH*GAU*(1.16e-008*sky130_fd_pr__nfet_05v0_nvt__toxe_mult*(sky130_fd_pr__nfet_05v0_nvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__nfet_05v0_nvt__rshn_mult'
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__esd_nfet_05v0_nvt__vth0_slope_spectre)
+ vth0 = '0.06+sky130_fd_pr__nfet_05v0_nvt__vth0_diff_1+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_05v0_nvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.364
+ k2 = '0.043475+sky130_fd_pr__nfet_05v0_nvt__k2_diff_1'
+ k3 = 1.4
+ dvt0 = 5.7
+ dvt1 = 0.21851
+ dvt2 = 0.04
+ dvt0w = 7.7
+ dvt1w = 1272000.0
+ dvt2w = -0.032
+ w0 = 0.0
+ k3b = -0.58
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = -1.2362266e-14
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '73076+sky130_fd_pr__nfet_05v0_nvt__vsat_diff_1'
+ ua = '8.4094e-010+sky130_fd_pr__nfet_05v0_nvt__ua_diff_1'
+ ub = '1.2348e-018+sky130_fd_pr__nfet_05v0_nvt__ub_diff_1'
+ uc = 2.9976e-11
+ rdsw = '430+sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_1'
+ prwb = 0.0
+ prwg = 1.0e-12
+ wr = 1.0
+ u0 = '0.049769+sky130_fd_pr__nfet_05v0_nvt__u0_diff_1'
+ a0 = '0.0832+sky130_fd_pr__nfet_05v0_nvt__a0_diff_1'
+ keta = '-0.019904+sky130_fd_pr__nfet_05v0_nvt__keta_diff_1'
+ a1 = 0.0
+ a2 = 0.96293372
+ ags = '0.70396+sky130_fd_pr__nfet_05v0_nvt__ags_diff_1'
+ b0 = '3.3993e-007+sky130_fd_pr__nfet_05v0_nvt__b0_diff_1'
+ b1 = '0+sky130_fd_pr__nfet_05v0_nvt__b1_diff_1'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__esd_nfet_05v0_nvt__voff_slope_spectre)
+ voff = '0+sky130_fd_pr__nfet_05v0_nvt__voff_diff_1+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_05v0_nvt__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__esd_nfet_05v0_nvt__nfactor_slope_spectre)
+ nfactor = '0.63313+sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_1+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_05v0_nvt__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = '0+sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_1'
+ cit = 9.2584123e-8
+ cdsc = 0.0
+ cdscb = 1.4150948e-7
+ cdscd = 1.5e-5
+ eta0 = '9+sky130_fd_pr__nfet_05v0_nvt__eta0_diff_1'
+ etab = -0.00021692
+ dsub = 0.42
* BSIM4 - Sub-threshold parameters
+ voffl = 1.9445332e-8
+ minv = 0.0
* Rout Parameters
+ pclm = '0.11748+sky130_fd_pr__nfet_05v0_nvt__pclm_diff_1'
+ pdiblc1 = 8.833e-7
+ pdiblc2 = 0.0002
+ pdiblcb = 0.0
+ drout = 0.13139
+ pscbe1 = 2.4476e+8
+ pscbe2 = 3.84e-9
+ pvag = 4.5419436
+ delta = 0.007
+ alpha0 = 2.01e-6
+ alpha1 = 0.093632
+ beta0 = 19.448
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0.0068+sky130_fd_pr__nfet_05v0_nvt__pdits_diff_1'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_1'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = '-0.35858+sky130_fd_pr__nfet_05v0_nvt__kt1_diff_1'
+ kt2 = -0.016016
+ at = 22800.0
+ ute = -1.7861
+ ua1 = 4.4e-10
+ ub1 = -1.6252e-18
+ uc1 = -3.94e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.5764
+ jss = 0.00042966
+ jsws = 8.040000000000001e-10
+ xtis = 0.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019685
+ tpbsw = 0.001
+ tpbswg = 0.0
+ tcj = 0.00083
+ tcjsw = 0.0
+ tcjswg = 0.0
+ cgdo = '3.473e-010*sky130_fd_pr__nfet_05v0_nvt__overlap_mult'
+ cgso = '3.473e-010*sky130_fd_pr__nfet_05v0_nvt__overlap_mult'
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '5e-011*sky130_fd_pr__nfet_05v0_nvt__overlap_mult'
+ cgdl = '5e-011*sky130_fd_pr__nfet_05v0_nvt__overlap_mult'
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = '7.6493e-008+sky130_fd_pr__nfet_05v0_nvt__dlc_diff+sky130_fd_pr__nfet_05v0_nvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__nfet_05v0_nvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 1.16
+ moin = 15.0
+ noff = 4.0
+ voffcv = 0.216
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.0008602*sky130_fd_pr__nfet_05v0_nvt__ajunction_mult'
+ mjs = 0.28329
+ pbs = 0.66345
+ cjsws = '8.5152e-011*sky130_fd_pr__nfet_05v0_nvt__pjunction_mult'
+ mjsws = 0.057926
+ pbsws = 1.0
+ cjswgs = '3.58e-011*sky130_fd_pr__nfet_05v0_nvt__pjunction_mult'
+ mjswgs = 0.33
+ pbswgs = 0.2442
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__nfet_05v0_nvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__nfet_05v0_nvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__nfet_05v0_nvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__nfet_05v0_nvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__nfet_05v0_nvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__nfet_05v0_nvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__nfet_05v0_nvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__nfet_05v0_nvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__esd_nfet_05v0_nvt__model.2 nmos
* DC IV MOS Parameters
+ lmin = 8.95e-07 lmax = 9.05e-07 wmin = 9.995e-06 wmax = 1.0005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '6.93e-008+sky130_fd_pr__nfet_05v0_nvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '4.5e-008+sky130_fd_pr__nfet_05v0_nvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.6e-9
+ dwb = 1.92e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.8
+ rnoib = 0.38
+ tnoia = 7.6e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__esd_nfet_05v0_nvt__toxe_slope_spectre)
+ toxe = '1.16e-008*sky130_fd_pr__nfet_05v0_nvt__toxe_mult+MC_MM_SWITCH*GAU*(1.16e-008*sky130_fd_pr__nfet_05v0_nvt__toxe_mult*(sky130_fd_pr__nfet_05v0_nvt__toxe_slope2/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__nfet_05v0_nvt__rshn_mult'
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__esd_nfet_05v0_nvt__vth0_slope_spectre)
+ vth0 = '0.062+sky130_fd_pr__nfet_05v0_nvt__vth0_diff_2+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_05v0_nvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.364
+ k2 = '0.038817+sky130_fd_pr__nfet_05v0_nvt__k2_diff_2'
+ k3 = 1.4
+ dvt0 = 5.7
+ dvt1 = 0.21851
+ dvt2 = 0.04
+ dvt0w = 7.7
+ dvt1w = 1272000.0
+ dvt2w = -0.032
+ w0 = 0.0
+ k3b = -0.58
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = -1.2362266e-14
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '74500+sky130_fd_pr__nfet_05v0_nvt__vsat_diff_2'
+ ua = '9.1406e-010+sky130_fd_pr__nfet_05v0_nvt__ua_diff_2'
+ ub = '1.2863e-018+sky130_fd_pr__nfet_05v0_nvt__ub_diff_2'
+ uc = 3.2583e-11
+ rdsw = '430+sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_2'
+ prwb = 0.0
+ prwg = 1.0e-12
+ wr = 1.0
+ u0 = '0.050801+sky130_fd_pr__nfet_05v0_nvt__u0_diff_2'
+ a0 = '0.08+sky130_fd_pr__nfet_05v0_nvt__a0_diff_2'
+ keta = '-0.019904+sky130_fd_pr__nfet_05v0_nvt__keta_diff_2'
+ a1 = 0.0
+ a2 = 0.96293372
+ ags = '0.87995+sky130_fd_pr__nfet_05v0_nvt__ags_diff_2'
+ b0 = '3.3993e-007+sky130_fd_pr__nfet_05v0_nvt__b0_diff_2'
+ b1 = '0+sky130_fd_pr__nfet_05v0_nvt__b1_diff_2'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__esd_nfet_05v0_nvt__voff_slope_spectre)
+ voff = '0+sky130_fd_pr__nfet_05v0_nvt__voff_diff_2+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_05v0_nvt__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__esd_nfet_05v0_nvt__nfactor_slope_spectre)
+ nfactor = '0.63313+sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_2+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_05v0_nvt__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = '0+sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_2'
+ cit = 9.2584123e-8
+ cdsc = 0.0
+ cdscb = 1.4150948e-7
+ cdscd = 1.5e-5
+ eta0 = '9+sky130_fd_pr__nfet_05v0_nvt__eta0_diff_2'
+ etab = -0.00021692
+ dsub = 0.42
* BSIM4 - Sub-threshold parameters
+ voffl = 1.9445332e-8
+ minv = 0.0
* Rout Parameters
+ pclm = '0.11748+sky130_fd_pr__nfet_05v0_nvt__pclm_diff_2'
+ pdiblc1 = 8.833e-7
+ pdiblc2 = 0.0002
+ pdiblcb = 0.0
+ drout = 0.13139
+ pscbe1 = 2.4476e+8
+ pscbe2 = 3.84e-9
+ pvag = 4.5419436
+ delta = 0.007
+ alpha0 = 2.1079e-6
+ alpha1 = 0.1232
+ beta0 = 25.668
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0.0002+sky130_fd_pr__nfet_05v0_nvt__pdits_diff_2'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_2'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = '-0.37322+sky130_fd_pr__nfet_05v0_nvt__kt1_diff_2'
+ kt2 = -0.01144
+ at = 19488.0
+ ute = -1.464
+ ua1 = 1.0e-9
+ ub1 = -7.128e-19
+ uc1 = 1.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.5764
+ jss = 0.00042966
+ jsws = 8.040000000000001e-10
+ xtis = 0.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019685
+ tpbsw = 0.001
+ tpbswg = 0.0
+ tcj = 0.00083
+ tcjsw = 0.0
+ tcjswg = 0.0
+ cgdo = '3.473e-010*sky130_fd_pr__nfet_05v0_nvt__overlap_mult'
+ cgso = '3.473e-010*sky130_fd_pr__nfet_05v0_nvt__overlap_mult'
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '5e-011*sky130_fd_pr__nfet_05v0_nvt__overlap_mult'
+ cgdl = '5e-011*sky130_fd_pr__nfet_05v0_nvt__overlap_mult'
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = '7.6493e-008+sky130_fd_pr__nfet_05v0_nvt__dlc_diff+sky130_fd_pr__nfet_05v0_nvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__nfet_05v0_nvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 1.16
+ moin = 15.0
+ noff = 4.0
+ voffcv = 0.216
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.0008602*sky130_fd_pr__nfet_05v0_nvt__ajunction_mult'
+ mjs = 0.28329
+ pbs = 0.66345
+ cjsws = '8.5152e-011*sky130_fd_pr__nfet_05v0_nvt__pjunction_mult'
+ mjsws = 0.057926
+ pbsws = 1.0
+ cjswgs = '3.58e-011*sky130_fd_pr__nfet_05v0_nvt__pjunction_mult'
+ mjswgs = 0.33
+ pbswgs = 0.2442
* Stress Parameters
+ saref = 2.54e-6
+ sbref = 2.54e-6
+ wlod = '0+sky130_fd_pr__nfet_05v0_nvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__nfet_05v0_nvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__nfet_05v0_nvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__nfet_05v0_nvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__nfet_05v0_nvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__nfet_05v0_nvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__nfet_05v0_nvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__nfet_05v0_nvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__esd_nfet_05v0_nvt
