* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param GAU = AGAUSS(0,1.0,1)
.param sky130_fd_pr__special_nfet_01v8__toxe_slope_spectre = 0.0
.param sky130_fd_pr__special_nfet_01v8__vth0_slope_spectre = 0.0
.param sky130_fd_pr__special_nfet_01v8__voff_slope_spectre = 0.0
.param sky130_fd_pr__special_nfet_01v8__nfactor_slope_spectre = 0.0
* statistics '
*   process '
*   '
*   mismatch '
*     vary sky130_fd_pr__special_nfet_01v8__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_nfet_01v8__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_nfet_01v8__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_nfet_01v8__nfactor_slope_spectre dist=gauss std = 1.0
*   '
* '
.subckt  sky130_fd_pr__special_nfet_01v8 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__special_nfet_01v8 d g s b sky130_fd_pr__special_nfet_01v8__model l = 'l' w = 'w' nf = 'nf' ad = 'ad' as = 'as' pd = 'pd' ps = 'ps' nrd = 'nrd' nrs = 'nrs' sa = 'sa' sb = 'sb' sd = 'sd'
.model sky130_fd_pr__special_nfet_01v8__model.0 nmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 3.59e-07 wmax = 3.61e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__special_nfet_01v8__toxe_slope_spectre)
+ toxe = '4.148e-09*sky130_fd_pr__special_nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__special_nfet_01v8__toxe_mult*(sky130_fd_pr__special_nfet_01v8__toxe_slope/sqrt(l*w*mult)))'
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = '1.0*sky130_fd_pr__special_nfet_01v8__rshn_mult'
+ rshg = 0.1
* Basic Model Parameters
+ wint = '2.1859e-08+sky130_fd_pr__special_nfet_01v8__wint_diff'
+ lint = '1.1932e-08+sky130_fd_pr__special_nfet_01v8__lint_diff'
*(mismatch parameter sky130_fd_pr__special_nfet_01v8__vth0_slope_spectre)
+ vth0 = '0.294216+sky130_fd_pr__special_nfet_01v8__vth0_diff_0+MC_MM_SWITCH*GAU*(sky130_fd_pr__special_nfet_01v8__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.90707349
+ k2 = '-0.164979+sky130_fd_pr__special_nfet_01v8__k2_diff_0'
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.745709255106775
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__special_nfet_01v8__voff_slope_spectre)
+ voff = '-0.20753+sky130_fd_pr__special_nfet_01v8__voff_diff_0+MC_MM_SWITCH*GAU*(sky130_fd_pr__special_nfet_01v8__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.11251750684601+sky130_fd_pr__special_nfet_01v8__nfactor_diff_0'
+ eta0 = '0.0+sky130_fd_pr__special_nfet_01v8__eta0_diff_0'
+ etab = -0.043998
+ u0 = '0.0420786+sky130_fd_pr__special_nfet_01v8__u0_diff_0'
+ ua = '-1.21575137545398e-09+sky130_fd_pr__special_nfet_01v8__ua_diff_0'
+ ub = '3.09344567610299e-18+sky130_fd_pr__special_nfet_01v8__ub_diff_0'
+ uc = 5.40303933016111e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = '205055.7+sky130_fd_pr__special_nfet_01v8__vsat_diff_0'
+ a0 = '1.5+sky130_fd_pr__special_nfet_01v8__a0_diff_0'
+ ags = '1.25+sky130_fd_pr__special_nfet_01v8__ags_diff_0'
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = '0.0+sky130_fd_pr__special_nfet_01v8__b0_diff_0'
+ b1 = '0.0+sky130_fd_pr__special_nfet_01v8__b1_diff_0'
+ keta = '-0.140717411247685+sky130_fd_pr__special_nfet_01v8__keta_diff_0'
+ dwg = 0.0
+ dwb = 0.0
+ pclm = '0.129289552416565+sky130_fd_pr__special_nfet_01v8__pclm_diff_0'
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = '0.0+sky130_fd_pr__special_nfet_01v8__pdits_diff_0'
+ pditsl = 0.0
+ pditsd = '0.0+sky130_fd_pr__special_nfet_01v8__pditsd_diff_0'
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = '65.968+sky130_fd_pr__special_nfet_01v8__rdsw_diff_0'
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.99999998238709e-8
+ alpha1 = 0.85
+ beta0 = 13.8499999988778
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = '1.0494e-08+sky130_fd_pr__special_nfet_01v8__dlc_diff+sky130_fd_pr__special_nfet_01v8__dlc_rotweak'
+ dwc = '0.0+sky130_fd_pr__special_nfet_01v8__dwc_diff'
+ xpart = 0.0
+ cgso = '2.54e-10*sky130_fd_pr__special_nfet_01v8__overlap_mult'
+ cgdo = '2.54e-10*sky130_fd_pr__special_nfet_01v8__overlap_mult'
+ cgbo = 1.0e-13
+ cgdl = '0.0*sky130_fd_pr__special_nfet_01v8__overlap_mult'
+ cgsl = '0.0*sky130_fd_pr__special_nfet_01v8__overlap_mult'
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = '0.0013459*sky130_fd_pr__special_nfet_01v8__ajunction_mult'
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = '3.6001e-11*sky130_fd_pr__special_nfet_01v8__pjunction_mult'
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = '2.3347e-10*sky130_fd_pr__special_nfet_01v8__pjunction_mult'
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = '-0.240960739938925+sky130_fd_pr__special_nfet_01v8__kt1_diff_0'
+ kt2 = -0.028878939
+ at = 53720.4870195945
+ ute = -1.19244645977108
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = '0.0+sky130_fd_pr__special_nfet_01v8__tvoff_diff_0'
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__special_nfet_01v8__model.0 nmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 3.89e-07 wmax = 3.91e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__special_nfet_01v8__toxe_slope_spectre)
+ toxe = '4.148e-09*sky130_fd_pr__special_nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__special_nfet_01v8__toxe_mult*(sky130_fd_pr__special_nfet_01v8__toxe_slope/sqrt(l*w*mult)))'
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = '1.0*sky130_fd_pr__special_nfet_01v8__rshn_mult'
+ rshg = 0.1
* Basic Model Parameters
+ wint = '2.1859e-08+sky130_fd_pr__special_nfet_01v8__wint_diff'
+ lint = '1.1932e-08+sky130_fd_pr__special_nfet_01v8__lint_diff'
*(mismatch parameter sky130_fd_pr__special_nfet_01v8__vth0_slope_spectre)
+ vth0 = '0.3288413+sky130_fd_pr__special_nfet_01v8__vth0_diff_1+MC_MM_SWITCH*GAU*(sky130_fd_pr__special_nfet_01v8__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.90707349
+ k2 = '-0.157868+sky130_fd_pr__special_nfet_01v8__k2_diff_1'
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.679435816074994
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__special_nfet_01v8__voff_slope_spectre)
+ voff = '-0.20753+sky130_fd_pr__special_nfet_01v8__voff_diff_1+MC_MM_SWITCH*GAU*(sky130_fd_pr__special_nfet_01v8__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.23668316177219+sky130_fd_pr__special_nfet_01v8__nfactor_diff_1'
+ eta0 = '0.0+sky130_fd_pr__special_nfet_01v8__eta0_diff_1'
+ etab = -0.043998
+ u0 = '0.0392402+sky130_fd_pr__special_nfet_01v8__u0_diff_1'
+ ua = '-1.20664055548599e-09+sky130_fd_pr__special_nfet_01v8__ua_diff_1'
+ ub = '2.8992935911323e-18+sky130_fd_pr__special_nfet_01v8__ub_diff_1'
+ uc = 6.17577815560697e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = '200231.2+sky130_fd_pr__special_nfet_01v8__vsat_diff_1'
+ a0 = '1.5+sky130_fd_pr__special_nfet_01v8__a0_diff_1'
+ ags = '1.25+sky130_fd_pr__special_nfet_01v8__ags_diff_1'
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = '0.0+sky130_fd_pr__special_nfet_01v8__b0_diff_1'
+ b1 = '0.0+sky130_fd_pr__special_nfet_01v8__b1_diff_1'
+ keta = '-0.114465726035654+sky130_fd_pr__special_nfet_01v8__keta_diff_1'
+ dwg = 0.0
+ dwb = 0.0
+ pclm = '0.137157029957607+sky130_fd_pr__special_nfet_01v8__pclm_diff_1'
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = '0.0+sky130_fd_pr__special_nfet_01v8__pdits_diff_1'
+ pditsl = 0.0
+ pditsd = '0.0+sky130_fd_pr__special_nfet_01v8__pditsd_diff_1'
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = '65.968+sky130_fd_pr__special_nfet_01v8__rdsw_diff_1'
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.99999998381496e-8
+ alpha1 = 0.85
+ beta0 = 13.8499999988803
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = '1.0494e-08+sky130_fd_pr__special_nfet_01v8__dlc_diff+sky130_fd_pr__special_nfet_01v8__dlc_rotweak'
+ dwc = '0.0+sky130_fd_pr__special_nfet_01v8__dwc_diff'
+ xpart = 0.0
+ cgso = '2.54e-10*sky130_fd_pr__special_nfet_01v8__overlap_mult'
+ cgdo = '2.54e-10*sky130_fd_pr__special_nfet_01v8__overlap_mult'
+ cgbo = 1.0e-13
+ cgdl = '0.0*sky130_fd_pr__special_nfet_01v8__overlap_mult'
+ cgsl = '0.0*sky130_fd_pr__special_nfet_01v8__overlap_mult'
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = '0.0013459*sky130_fd_pr__special_nfet_01v8__ajunction_mult'
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = '3.6001e-11*sky130_fd_pr__special_nfet_01v8__pjunction_mult'
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = '2.3347e-10*sky130_fd_pr__special_nfet_01v8__pjunction_mult'
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = '-0.240960739944239+sky130_fd_pr__special_nfet_01v8__kt1_diff_1'
+ kt2 = -0.028878939
+ at = 53720.4870179085
+ ute = -1.20689692868465
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = '0.0+sky130_fd_pr__special_nfet_01v8__tvoff_diff_1'
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.ends sky130_fd_pr__special_nfet_01v8
