* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param GAU = AGAUSS(0,1.0,1)
.param sky130_fd_pr__nfet_01v8__toxe_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__vth0_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__voff_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_01v8__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
* "special" standard cell nFET (w < 0.42um) is defined as a regular nFET because its model bins exist there.
.subckt  sky130_fd_pr__special_nfet_01v8 d g s b
+
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
xsky130_fd_pr__nfet_01v8 d g s b sky130_fd_pr__nfet_01v8 l = 'l' w = 'w' nf = 'nf' ad = 'ad' as = 'as' pd = 'pd' ps = 'ps' nrd = 'nrd' nrs = 'nrs' sa = 'sa' sb = 'sb' sd = 'sd'
.ends

.subckt  sky130_fd_pr__nfet_01v8 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__nfet_01v8 d g s b sky130_fd_pr__nfet_01v8__model l = 'l' w = 'w' nf = 'nf' ad = 'ad' as = 'as' pd = 'pd' ps = 'ps' nrd = 'nrd' nrs = 'nrs' sa = 'sa' sb = 'sb' sd = 'sd'
.model sky130_fd_pr__nfet_01v8__model.0 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.255e-06 wmax = 1.265e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.49439+sky130_fd_pr__nfet_01v8__vth0_diff_0+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.12949+sky130_fd_pr__nfet_01v8__k2_diff_0}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {176320+sky130_fd_pr__nfet_01v8__vsat_diff_0}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_0}
+ ub = {2.1846e-018+sky130_fd_pr__nfet_01v8__ub_diff_0}
+ uc = 8.1022e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_0}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.030197+sky130_fd_pr__nfet_01v8__u0_diff_0}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_0}
+ keta = {0+sky130_fd_pr__nfet_01v8__keta_diff_0}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_0}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_0}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_0}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_0+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {2.015+sky130_fd_pr__nfet_01v8__nfactor_diff_0+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_0}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0.00069413878+sky130_fd_pr__nfet_01v8__eta0_diff_0}
+ etab = -0.043998
+ dsub = 0.45862506
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.14094+sky130_fd_pr__nfet_01v8__pclm_diff_0}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.85
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_0}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_0}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.22096074+sky130_fd_pr__nfet_01v8__kt1_diff_0}
+ kt2 = -0.028878939
+ at = 40720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.1 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.675e-06 wmax = 1.685e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.45777+sky130_fd_pr__nfet_01v8__vth0_diff_1+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.13489+sky130_fd_pr__nfet_01v8__k2_diff_1}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {176320+sky130_fd_pr__nfet_01v8__vsat_diff_1}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_1}
+ ub = {2.1006e-018+sky130_fd_pr__nfet_01v8__ub_diff_1}
+ uc = 6.4303e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_1}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.030197+sky130_fd_pr__nfet_01v8__u0_diff_1}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_1}
+ keta = {0+sky130_fd_pr__nfet_01v8__keta_diff_1}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_1}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_1}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_1}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_1+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {2.015+sky130_fd_pr__nfet_01v8__nfactor_diff_1+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_1}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0.00069413878+sky130_fd_pr__nfet_01v8__eta0_diff_1}
+ etab = -0.043998
+ dsub = 0.45862506
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.14094+sky130_fd_pr__nfet_01v8__pclm_diff_1}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.82
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_1}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_1}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.22096074+sky130_fd_pr__nfet_01v8__kt1_diff_1}
+ kt2 = -0.028878939
+ at = 60720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.2 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.57666+sky130_fd_pr__nfet_01v8__vth0_diff_2+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47926744
+ k2 = {-0.00734+sky130_fd_pr__nfet_01v8__k2_diff_2}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {90000+sky130_fd_pr__nfet_01v8__vsat_diff_2}
+ ua = {-1.3915e-009+sky130_fd_pr__nfet_01v8__ua_diff_2}
+ ub = {1.9256e-018+sky130_fd_pr__nfet_01v8__ub_diff_2}
+ uc = 7.0144e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_2}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.024597+sky130_fd_pr__nfet_01v8__u0_diff_2}
+ a0 = {0.4182+sky130_fd_pr__nfet_01v8__a0_diff_2}
+ keta = {0.0095396+sky130_fd_pr__nfet_01v8__keta_diff_2}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.72513+sky130_fd_pr__nfet_01v8__ags_diff_2}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_2}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_2}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.15134+sky130_fd_pr__nfet_01v8__voff_diff_2+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {0.84726+sky130_fd_pr__nfet_01v8__nfactor_diff_2+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_2}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.0025313+sky130_fd_pr__nfet_01v8__eta0_diff_2}
+ etab = -0.084375
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.68831+sky130_fd_pr__nfet_01v8__pclm_diff_2}
+ pdiblc1 = 0.33870462
+ pdiblc2 = 0.005806679
+ pdiblcb = -0.04937254
+ drout = 0.39729981
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.88e-8
+ alpha1 = 0.697
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_2}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_2}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25664+sky130_fd_pr__nfet_01v8__kt1_diff_2}
+ kt2 = -0.036226822
+ at = 85715.0
+ ute = -1.0468
+ ua1 = 1.2463e-9
+ ub1 = -7.6772e-19
+ uc1 = 1.8046812e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.3 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.55639+sky130_fd_pr__nfet_01v8__vth0_diff_3+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53942222
+ k2 = {-0.02714132+sky130_fd_pr__nfet_01v8__k2_diff_3}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_3}
+ ua = {-1.1570455e-009+sky130_fd_pr__nfet_01v8__ua_diff_3}
+ ub = {1.8354e-018+sky130_fd_pr__nfet_01v8__ub_diff_3}
+ uc = 5.4094e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_3}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.02701+sky130_fd_pr__nfet_01v8__u0_diff_3}
+ a0 = {1.008+sky130_fd_pr__nfet_01v8__a0_diff_3}
+ keta = {-0.0088430972+sky130_fd_pr__nfet_01v8__keta_diff_3}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.50628+sky130_fd_pr__nfet_01v8__ags_diff_3}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_3}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_3}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.12584821+sky130_fd_pr__nfet_01v8__voff_diff_3+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.5798554+sky130_fd_pr__nfet_01v8__nfactor_diff_3+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_3}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_3}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.55709+sky130_fd_pr__nfet_01v8__pclm_diff_3}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0052969163
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_3}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_3}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.29168+sky130_fd_pr__nfet_01v8__kt1_diff_3}
+ kt2 = -0.017698782
+ at = 111200.0
+ ute = -0.42247
+ ua1 = 3.6107e-9
+ ub1 = -2.7362e-18
+ uc1 = -3.0219439e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.4 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.54021+sky130_fd_pr__nfet_01v8__vth0_diff_4+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.49025322
+ k2 = {-0.012213166+sky130_fd_pr__nfet_01v8__k2_diff_4}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_4}
+ ua = {-7.0340514e-010+sky130_fd_pr__nfet_01v8__ua_diff_4}
+ ub = {1.391e-018+sky130_fd_pr__nfet_01v8__ub_diff_4}
+ uc = 2.5377e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_4}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.02967+sky130_fd_pr__nfet_01v8__u0_diff_4}
+ a0 = {1.2+sky130_fd_pr__nfet_01v8__a0_diff_4}
+ keta = {0.0097600722+sky130_fd_pr__nfet_01v8__keta_diff_4}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.3478+sky130_fd_pr__nfet_01v8__ags_diff_4}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_4}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_4}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.1060102+sky130_fd_pr__nfet_01v8__voff_diff_4+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_4+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_4}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_4}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.53316+sky130_fd_pr__nfet_01v8__pclm_diff_4}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0033446417
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.452285e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_4}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_4}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.29371+sky130_fd_pr__nfet_01v8__kt1_diff_4}
+ kt2 = -0.020698378
+ at = 140000.0
+ ute = -1.0855
+ ua1 = 1.4555e-9
+ ub1 = -9.4827e-19
+ uc1 = -1.8284811e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.5 nmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.53654+sky130_fd_pr__nfet_01v8__vth0_diff_5+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47351598
+ k2 = {-0.0058110531+sky130_fd_pr__nfet_01v8__k2_diff_5}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_5}
+ ua = {-6.6692005e-010+sky130_fd_pr__nfet_01v8__ua_diff_5}
+ ub = {1.3895e-018+sky130_fd_pr__nfet_01v8__ub_diff_5}
+ uc = 2.5799e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_5}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.030717+sky130_fd_pr__nfet_01v8__u0_diff_5}
+ a0 = {1.32+sky130_fd_pr__nfet_01v8__a0_diff_5}
+ keta = {-0.0015333577+sky130_fd_pr__nfet_01v8__keta_diff_5}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.36348+sky130_fd_pr__nfet_01v8__ags_diff_5}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_5}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_5}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.11141737+sky130_fd_pr__nfet_01v8__voff_diff_5+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_5+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_5}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_5}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.083531+sky130_fd_pr__nfet_01v8__pclm_diff_5}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0031503727
+ pdiblcb = -2.2185512
+ drout = 0.56
+ pscbe1 = 7.615138e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_5}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_5}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.29248+sky130_fd_pr__nfet_01v8__kt1_diff_5}
+ kt2 = -0.020636654
+ at = 140000.0
+ ute = -1.2877
+ ua1 = 1.3536e-9
+ ub1 = -9.4206e-19
+ uc1 = -2.4408323e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.6 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.47461+sky130_fd_pr__nfet_01v8__vth0_diff_6+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.12949+sky130_fd_pr__nfet_01v8__k2_diff_6}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {183370+sky130_fd_pr__nfet_01v8__vsat_diff_6}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_6}
+ ub = {2.1846e-018+sky130_fd_pr__nfet_01v8__ub_diff_6}
+ uc = 8.1022e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_6}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.030197+sky130_fd_pr__nfet_01v8__u0_diff_6}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_6}
+ keta = {0+sky130_fd_pr__nfet_01v8__keta_diff_6}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_6}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_6}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_6}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_6+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {2.015+sky130_fd_pr__nfet_01v8__nfactor_diff_6+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_6}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0.00069413878+sky130_fd_pr__nfet_01v8__eta0_diff_6}
+ etab = -0.043998
+ dsub = 0.45862506
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.12966+sky130_fd_pr__nfet_01v8__pclm_diff_6}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.85
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_6}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_6}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.22096074+sky130_fd_pr__nfet_01v8__kt1_diff_6}
+ kt2 = -0.028878939
+ at = 40720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.7 nmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.50758+sky130_fd_pr__nfet_01v8__vth0_diff_7+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.13467+sky130_fd_pr__nfet_01v8__k2_diff_7}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {183370+sky130_fd_pr__nfet_01v8__vsat_diff_7}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_7}
+ ub = {2.1846e-018+sky130_fd_pr__nfet_01v8__ub_diff_7}
+ uc = 1.1019e-10
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_7}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.029997+sky130_fd_pr__nfet_01v8__u0_diff_7}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_7}
+ keta = {-0.039+sky130_fd_pr__nfet_01v8__keta_diff_7}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_7}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_7}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_7}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_7+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.209+sky130_fd_pr__nfet_01v8__nfactor_diff_7+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_7}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0.00069413878+sky130_fd_pr__nfet_01v8__eta0_diff_7}
+ etab = -0.043998
+ dsub = 0.45862506
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.12966+sky130_fd_pr__nfet_01v8__pclm_diff_7}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.16e-8
+ alpha1 = 0.85
+ beta0 = 14.08
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_7}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_7}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.24096074+sky130_fd_pr__nfet_01v8__kt1_diff_7}
+ kt2 = -0.028878939
+ at = 60720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.8 nmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.54308+sky130_fd_pr__nfet_01v8__vth0_diff_8+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.14006+sky130_fd_pr__nfet_01v8__k2_diff_8}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {175450+sky130_fd_pr__nfet_01v8__vsat_diff_8}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_8}
+ ub = {1.8655e-018+sky130_fd_pr__nfet_01v8__ub_diff_8}
+ uc = 9.256e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_8}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.030197+sky130_fd_pr__nfet_01v8__u0_diff_8}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_8}
+ keta = {-0.083148+sky130_fd_pr__nfet_01v8__keta_diff_8}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_8}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_8}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_8}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.17848+sky130_fd_pr__nfet_01v8__voff_diff_8+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.209+sky130_fd_pr__nfet_01v8__nfactor_diff_8+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_8}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0.00069414+sky130_fd_pr__nfet_01v8__eta0_diff_8}
+ etab = -0.043998
+ dsub = 0.45863
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23857+sky130_fd_pr__nfet_01v8__pclm_diff_8}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.16e-8
+ alpha1 = 0.85
+ beta0 = 14.32
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_8}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_8}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.24096074+sky130_fd_pr__nfet_01v8__kt1_diff_8}
+ kt2 = -0.028878939
+ at = 28720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.9 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.57726635+sky130_fd_pr__nfet_01v8__vth0_diff_9+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56348836
+ k2 = {-0.040381304+sky130_fd_pr__nfet_01v8__k2_diff_9}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {131360+sky130_fd_pr__nfet_01v8__vsat_diff_9}
+ ua = {-1.4916409e-009+sky130_fd_pr__nfet_01v8__ua_diff_9}
+ ub = {2.08e-018+sky130_fd_pr__nfet_01v8__ub_diff_9}
+ uc = 7.754e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_9}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.024638+sky130_fd_pr__nfet_01v8__u0_diff_9}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_9}
+ keta = {-0.031644245+sky130_fd_pr__nfet_01v8__keta_diff_9}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.0952+sky130_fd_pr__nfet_01v8__ags_diff_9}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_9}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_9}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.14543985+sky130_fd_pr__nfet_01v8__voff_diff_9+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.7093856+sky130_fd_pr__nfet_01v8__nfactor_diff_9+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_9}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.49+sky130_fd_pr__nfet_01v8__eta0_diff_9}
+ etab = -0.0003125
+ dsub = 0.31335602
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.5+sky130_fd_pr__nfet_01v8__pclm_diff_9}
+ pdiblc1 = 0.14211905
+ pdiblc2 = 0.0016058161
+ pdiblcb = -0.025
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_9}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_9}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27076249+sky130_fd_pr__nfet_01v8__kt1_diff_9}
+ kt2 = -0.036350227
+ at = 50130.388
+ ute = -1.2259453
+ ua1 = 1.0936141e-9
+ ub1 = -6.797397e-19
+ uc1 = 3.9201824e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.10 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.995e-06 wmax = 2.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.45777+sky130_fd_pr__nfet_01v8__vth0_diff_10+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.13489+sky130_fd_pr__nfet_01v8__k2_diff_10}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {173320+sky130_fd_pr__nfet_01v8__vsat_diff_10}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_10}
+ ub = {2.1881e-018+sky130_fd_pr__nfet_01v8__ub_diff_10}
+ uc = 8.244e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_10}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.030197+sky130_fd_pr__nfet_01v8__u0_diff_10}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_10}
+ keta = {0.018418+sky130_fd_pr__nfet_01v8__keta_diff_10}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_10}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_10}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_10}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_10+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {2.015+sky130_fd_pr__nfet_01v8__nfactor_diff_10+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_10}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0.00069413878+sky130_fd_pr__nfet_01v8__eta0_diff_10}
+ etab = -0.043998
+ dsub = 0.45862506
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.1532+sky130_fd_pr__nfet_01v8__pclm_diff_10}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_10}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_10}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.24096074+sky130_fd_pr__nfet_01v8__kt1_diff_10}
+ kt2 = -0.028878939
+ at = 60720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.11 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.56797+sky130_fd_pr__nfet_01v8__vth0_diff_11+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.50655102
+ k2 = {-0.017147679+sky130_fd_pr__nfet_01v8__k2_diff_11}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {75585+sky130_fd_pr__nfet_01v8__vsat_diff_11}
+ ua = {-1.4807062e-009+sky130_fd_pr__nfet_01v8__ua_diff_11}
+ ub = {2.189e-018+sky130_fd_pr__nfet_01v8__ub_diff_11}
+ uc = 7.4874e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_11}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.025492+sky130_fd_pr__nfet_01v8__u0_diff_11}
+ a0 = {0.93+sky130_fd_pr__nfet_01v8__a0_diff_11}
+ keta = {-0.051315+sky130_fd_pr__nfet_01v8__keta_diff_11}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.2+sky130_fd_pr__nfet_01v8__ags_diff_11}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_11}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_11}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.13377387+sky130_fd_pr__nfet_01v8__voff_diff_11+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.3879762+sky130_fd_pr__nfet_01v8__nfactor_diff_11+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_11}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.00253125+sky130_fd_pr__nfet_01v8__eta0_diff_11}
+ etab = -0.084375
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.88922+sky130_fd_pr__nfet_01v8__pclm_diff_11}
+ pdiblc1 = 0.62056999
+ pdiblc2 = 0.0032799909
+ pdiblcb = -0.0001916735
+ drout = 0.26
+ pscbe1 = 4.1970592e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.88e-8
+ alpha1 = 1.071
+ beta0 = 14.529
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_11}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_11}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25495+sky130_fd_pr__nfet_01v8__kt1_diff_11}
+ kt2 = -0.035831378
+ at = 65630.0
+ ute = -1.1735
+ ua1 = 1.6342407e-9
+ ub1 = -1.4490891e-18
+ uc1 = -1.5193288e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.12 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.54406+sky130_fd_pr__nfet_01v8__vth0_diff_12+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56914885
+ k2 = {-0.043416987+sky130_fd_pr__nfet_01v8__k2_diff_12}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_12}
+ ua = {-8.0325375e-010+sky130_fd_pr__nfet_01v8__ua_diff_12}
+ ub = {1.7925e-018+sky130_fd_pr__nfet_01v8__ub_diff_12}
+ uc = 6.411e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_12}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.032582+sky130_fd_pr__nfet_01v8__u0_diff_12}
+ a0 = {1.4904+sky130_fd_pr__nfet_01v8__a0_diff_12}
+ keta = {0.00038915367+sky130_fd_pr__nfet_01v8__keta_diff_12}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.69201+sky130_fd_pr__nfet_01v8__ags_diff_12}
+ b0 = {2.1073e-024+sky130_fd_pr__nfet_01v8__b0_diff_12}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_12}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.10092566+sky130_fd_pr__nfet_01v8__voff_diff_12+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_12+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_12}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_12}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.50406+sky130_fd_pr__nfet_01v8__pclm_diff_12}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0048489026
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.9166137e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_12}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_12}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.32212+sky130_fd_pr__nfet_01v8__kt1_diff_12}
+ kt2 = -0.041614362
+ at = 115100.0
+ ute = -1.5856
+ ua1 = 5.4706e-10
+ ub1 = -4.0777e-19
+ uc1 = 4.4867589e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.13 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.53706+sky130_fd_pr__nfet_01v8__vth0_diff_13+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55462267
+ k2 = {-0.037104101+sky130_fd_pr__nfet_01v8__k2_diff_13}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_13}
+ ua = {-6.6780205e-010+sky130_fd_pr__nfet_01v8__ua_diff_13}
+ ub = {1.6832e-018+sky130_fd_pr__nfet_01v8__ub_diff_13}
+ uc = 6.0646e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_13}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.033867+sky130_fd_pr__nfet_01v8__u0_diff_13}
+ a0 = {1.26+sky130_fd_pr__nfet_01v8__a0_diff_13}
+ keta = {-0.00068634+sky130_fd_pr__nfet_01v8__keta_diff_13}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.42318+sky130_fd_pr__nfet_01v8__ags_diff_13}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_13}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_13}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.10370521+sky130_fd_pr__nfet_01v8__voff_diff_13+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_13+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_13}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_13}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.48885+sky130_fd_pr__nfet_01v8__pclm_diff_13}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0034912054
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_13}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_13}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.31856+sky130_fd_pr__nfet_01v8__kt1_diff_13}
+ kt2 = -0.042161763
+ at = 140000.0
+ ute = -1.763
+ ua1 = 2.8663405e-10
+ ub1 = -3.5073801e-19
+ uc1 = 2.7151174e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.14 nmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.52903+sky130_fd_pr__nfet_01v8__vth0_diff_14+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55146741
+ k2 = {-0.034414452+sky130_fd_pr__nfet_01v8__k2_diff_14}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_14}
+ ua = {-7.1064448e-010+sky130_fd_pr__nfet_01v8__ua_diff_14}
+ ub = {1.7147e-018+sky130_fd_pr__nfet_01v8__ub_diff_14}
+ uc = 7.0972e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_14}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.033266+sky130_fd_pr__nfet_01v8__u0_diff_14}
+ a0 = {1.38+sky130_fd_pr__nfet_01v8__a0_diff_14}
+ keta = {-0.0056579+sky130_fd_pr__nfet_01v8__keta_diff_14}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.43785+sky130_fd_pr__nfet_01v8__ags_diff_14}
+ b0 = {2.1073e-024+sky130_fd_pr__nfet_01v8__b0_diff_14}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_14}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.10574827+sky130_fd_pr__nfet_01v8__voff_diff_14+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_14+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_14}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_14}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.083531+sky130_fd_pr__nfet_01v8__pclm_diff_14}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0024625373
+ pdiblcb = -2.5116166
+ drout = 0.56
+ pscbe1 = 7.9351578e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_14}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_14}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.31634+sky130_fd_pr__nfet_01v8__kt1_diff_14}
+ kt2 = -0.041061662
+ at = 140000.0
+ ute = -1.7903
+ ua1 = 3.3088e-10
+ ub1 = -4.2516e-19
+ uc1 = 1.5167332e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.15 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.45777+sky130_fd_pr__nfet_01v8__vth0_diff_15+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.14051+sky130_fd_pr__nfet_01v8__k2_diff_15}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {166650+sky130_fd_pr__nfet_01v8__vsat_diff_15}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_15}
+ ub = {2.2793e-018+sky130_fd_pr__nfet_01v8__ub_diff_15}
+ uc = 5.9739e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_15}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.030197+sky130_fd_pr__nfet_01v8__u0_diff_15}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_15}
+ keta = {0.018418+sky130_fd_pr__nfet_01v8__keta_diff_15}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_15}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_15}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_15}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.18204+sky130_fd_pr__nfet_01v8__voff_diff_15+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {2.2389+sky130_fd_pr__nfet_01v8__nfactor_diff_15+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_15}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0.00069413878+sky130_fd_pr__nfet_01v8__eta0_diff_15}
+ etab = -0.051161
+ dsub = 0.45862506
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.15958+sky130_fd_pr__nfet_01v8__pclm_diff_15}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_15}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_15}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25096074+sky130_fd_pr__nfet_01v8__kt1_diff_15}
+ kt2 = -0.028878939
+ at = 60720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.16 nmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.49439+sky130_fd_pr__nfet_01v8__vth0_diff_16+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.14051+sky130_fd_pr__nfet_01v8__k2_diff_16}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {153320+sky130_fd_pr__nfet_01v8__vsat_diff_16}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_16}
+ ub = {2.1881e-018+sky130_fd_pr__nfet_01v8__ub_diff_16}
+ uc = 5.9739e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_16}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.030197+sky130_fd_pr__nfet_01v8__u0_diff_16}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_16}
+ keta = {-0.050739+sky130_fd_pr__nfet_01v8__keta_diff_16}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_16}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_16}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_16}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.18204+sky130_fd_pr__nfet_01v8__voff_diff_16+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.7911+sky130_fd_pr__nfet_01v8__nfactor_diff_16+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_16}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0.00069414+sky130_fd_pr__nfet_01v8__eta0_diff_16}
+ etab = -0.051161
+ dsub = 0.45863
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.25533+sky130_fd_pr__nfet_01v8__pclm_diff_16}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 14.25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_16}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_16}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25096074+sky130_fd_pr__nfet_01v8__kt1_diff_16}
+ kt2 = -0.028878939
+ at = 75720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.17 nmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.54854+sky130_fd_pr__nfet_01v8__vth0_diff_17+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.77890192
+ k2 = {-0.09820953+sky130_fd_pr__nfet_01v8__k2_diff_17}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {153850+sky130_fd_pr__nfet_01v8__vsat_diff_17}
+ ua = {-2.0950794e-009+sky130_fd_pr__nfet_01v8__ua_diff_17}
+ ub = {2.3625e-018+sky130_fd_pr__nfet_01v8__ub_diff_17}
+ uc = 7.4412e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_17}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.0179+sky130_fd_pr__nfet_01v8__u0_diff_17}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_17}
+ keta = {-0.039919373+sky130_fd_pr__nfet_01v8__keta_diff_17}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.019531+sky130_fd_pr__nfet_01v8__ags_diff_17}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_17}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_17}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.1450501+sky130_fd_pr__nfet_01v8__voff_diff_17+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.6674737+sky130_fd_pr__nfet_01v8__nfactor_diff_17+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_17}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.49+sky130_fd_pr__nfet_01v8__eta0_diff_17}
+ etab = -0.000625
+ dsub = 0.5734777
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.32133+sky130_fd_pr__nfet_01v8__pclm_diff_17}
+ pdiblc1 = 0.15540287
+ pdiblc2 = 0.0025814363
+ pdiblcb = -0.225
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.3e-6
+ alpha1 = 0.85
+ beta0 = 19.127
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_17}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_17}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.24632158+sky130_fd_pr__nfet_01v8__kt1_diff_17}
+ kt2 = -0.017111219
+ at = 22692.407
+ ute = -0.28054438
+ ua1 = 2.3883282e-9
+ ub1 = -1.4441988e-18
+ uc1 = 5.0765509e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.18 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.58344+sky130_fd_pr__nfet_01v8__vth0_diff_18+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57718752
+ k2 = {-0.044213929+sky130_fd_pr__nfet_01v8__k2_diff_18}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {124150+sky130_fd_pr__nfet_01v8__vsat_diff_18}
+ ua = {-1.5972244e-009+sky130_fd_pr__nfet_01v8__ua_diff_18}
+ ub = {2.14e-018+sky130_fd_pr__nfet_01v8__ub_diff_18}
+ uc = 7.5805e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_18}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.02368+sky130_fd_pr__nfet_01v8__u0_diff_18}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_18}
+ keta = {-0.035567981+sky130_fd_pr__nfet_01v8__keta_diff_18}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.1844+sky130_fd_pr__nfet_01v8__ags_diff_18}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_18}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_18}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.1394277+sky130_fd_pr__nfet_01v8__voff_diff_18+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8160129+sky130_fd_pr__nfet_01v8__nfactor_diff_18+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_18}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.49+sky130_fd_pr__nfet_01v8__eta0_diff_18}
+ etab = -0.000625
+ dsub = 0.32987125
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.4+sky130_fd_pr__nfet_01v8__pclm_diff_18}
+ pdiblc1 = 0.5
+ pdiblc2 = 0.0010936016
+ pdiblcb = -0.025
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.24e-6
+ alpha1 = 0.85
+ beta0 = 18.018
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_18}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_18}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27918368+sky130_fd_pr__nfet_01v8__kt1_diff_18}
+ kt2 = -0.03692268
+ at = 46593.516
+ ute = -1.2530532
+ ua1 = 1.0416734e-9
+ ub1 = -5.790873e-19
+ uc1 = 5.2032528e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.19 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.5565+sky130_fd_pr__nfet_01v8__vth0_diff_19+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57126962
+ k2 = {-0.046981026+sky130_fd_pr__nfet_01v8__k2_diff_19}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {83868+sky130_fd_pr__nfet_01v8__vsat_diff_19}
+ ua = {-1.4195372e-009+sky130_fd_pr__nfet_01v8__ua_diff_19}
+ ub = {2.14e-018+sky130_fd_pr__nfet_01v8__ub_diff_19}
+ uc = 5.0555e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_19}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.026261+sky130_fd_pr__nfet_01v8__u0_diff_19}
+ a0 = {1.38+sky130_fd_pr__nfet_01v8__a0_diff_19}
+ keta = {-0.066895435+sky130_fd_pr__nfet_01v8__keta_diff_19}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_19}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_19}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_19}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.12341816+sky130_fd_pr__nfet_01v8__voff_diff_19+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.6787831+sky130_fd_pr__nfet_01v8__nfactor_diff_19+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_19}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.00049393699+sky130_fd_pr__nfet_01v8__eta0_diff_19}
+ etab = -0.00042636116
+ dsub = 0.6209372
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.33434+sky130_fd_pr__nfet_01v8__pclm_diff_19}
+ pdiblc1 = 0.59602251
+ pdiblc2 = 0.0050495029
+ pdiblcb = -9.6868067e-5
+ drout = 0.26
+ pscbe1 = 6.7482021e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.84e-6
+ alpha1 = 0.884
+ beta0 = 16.909
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_19}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_19}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27358333+sky130_fd_pr__nfet_01v8__kt1_diff_19}
+ kt2 = -0.026425531
+ at = 62107.214
+ ute = -0.84493977
+ ua1 = 2.2952124e-9
+ ub1 = -1.5373115e-18
+ uc1 = 5.0612086e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.20 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.54545+sky130_fd_pr__nfet_01v8__vth0_diff_20+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56069487
+ k2 = {-0.041367273+sky130_fd_pr__nfet_01v8__k2_diff_20}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_20}
+ ua = {-8.2159816e-010+sky130_fd_pr__nfet_01v8__ua_diff_20}
+ ub = {1.9408e-018+sky130_fd_pr__nfet_01v8__ub_diff_20}
+ uc = 7.1836e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_20}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.034119+sky130_fd_pr__nfet_01v8__u0_diff_20}
+ a0 = {1.1616+sky130_fd_pr__nfet_01v8__a0_diff_20}
+ keta = {0.0013859955+sky130_fd_pr__nfet_01v8__keta_diff_20}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.59557+sky130_fd_pr__nfet_01v8__ags_diff_20}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_20}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_20}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.0991204+sky130_fd_pr__nfet_01v8__voff_diff_20+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_20+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_20}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.0005+sky130_fd_pr__nfet_01v8__eta0_diff_20}
+ etab = -0.00050000011
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.45442+sky130_fd_pr__nfet_01v8__pclm_diff_20}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0050760312
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_20}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_20}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.3273+sky130_fd_pr__nfet_01v8__kt1_diff_20}
+ kt2 = -0.042188396
+ at = 116170.0
+ ute = -1.6863
+ ua1 = 4.6161e-10
+ ub1 = -4.6448e-19
+ uc1 = 3.5002802e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.21 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.53656+sky130_fd_pr__nfet_01v8__vth0_diff_21+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55023127
+ k2 = {-0.035260333+sky130_fd_pr__nfet_01v8__k2_diff_21}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_21}
+ ua = {-7.3862315e-010+sky130_fd_pr__nfet_01v8__ua_diff_21}
+ ub = {1.8657e-018+sky130_fd_pr__nfet_01v8__ub_diff_21}
+ uc = 8.6636e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_21}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.034369+sky130_fd_pr__nfet_01v8__u0_diff_21}
+ a0 = {1.3104+sky130_fd_pr__nfet_01v8__a0_diff_21}
+ keta = {-0.0020009+sky130_fd_pr__nfet_01v8__keta_diff_21}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.51228+sky130_fd_pr__nfet_01v8__ags_diff_21}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_21}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_21}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.10282899+sky130_fd_pr__nfet_01v8__voff_diff_21+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_21+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_21}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_21}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.49027+sky130_fd_pr__nfet_01v8__pclm_diff_21}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0032336046
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.9893128e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_21}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_21}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.31714+sky130_fd_pr__nfet_01v8__kt1_diff_21}
+ kt2 = -0.041937248
+ at = 140000.0
+ ute = -1.7286
+ ua1 = 4.9161e-10
+ ub1 = -6.24e-19
+ uc1 = 2.0933495e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.22 nmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.52276+sky130_fd_pr__nfet_01v8__vth0_diff_22+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.54240333
+ k2 = {-0.031837301+sky130_fd_pr__nfet_01v8__k2_diff_22}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_22}
+ ua = {-7.2655782e-010+sky130_fd_pr__nfet_01v8__ua_diff_22}
+ ub = {1.6776e-018+sky130_fd_pr__nfet_01v8__ub_diff_22}
+ uc = 4.6783e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_22}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.033068+sky130_fd_pr__nfet_01v8__u0_diff_22}
+ a0 = {1.35+sky130_fd_pr__nfet_01v8__a0_diff_22}
+ keta = {-0.0061869508+sky130_fd_pr__nfet_01v8__keta_diff_22}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.39376+sky130_fd_pr__nfet_01v8__ags_diff_22}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_22}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_22}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.10408056+sky130_fd_pr__nfet_01v8__voff_diff_22+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_22+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_22}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_22}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.076882+sky130_fd_pr__nfet_01v8__pclm_diff_22}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0031936889
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.945303e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_22}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_22}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.3244+sky130_fd_pr__nfet_01v8__kt1_diff_22}
+ kt2 = -0.045509503
+ at = 140000.0
+ ute = -1.8837
+ ua1 = 2.591e-10
+ ub1 = -4.9785e-19
+ uc1 = 1.7026927e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.23 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.42361+sky130_fd_pr__nfet_01v8__vth0_diff_23+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90167256
+ k2 = {-0.12414+sky130_fd_pr__nfet_01v8__k2_diff_23}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {159280+sky130_fd_pr__nfet_01v8__vsat_diff_23}
+ ua = {-2.378e-009+sky130_fd_pr__nfet_01v8__ua_diff_23}
+ ub = {2.6241e-018+sky130_fd_pr__nfet_01v8__ub_diff_23}
+ uc = 4.1671e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_23}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.014112+sky130_fd_pr__nfet_01v8__u0_diff_23}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_23}
+ keta = {-0.059018+sky130_fd_pr__nfet_01v8__keta_diff_23}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_23}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_23}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_23}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.16464+sky130_fd_pr__nfet_01v8__voff_diff_23+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.9738+sky130_fd_pr__nfet_01v8__nfactor_diff_23+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_23}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.003456
+ eta0 = {0.00071353727+sky130_fd_pr__nfet_01v8__eta0_diff_23}
+ etab = -0.03833
+ dsub = 0.39261382
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.14349+sky130_fd_pr__nfet_01v8__pclm_diff_23}
+ pdiblc1 = 0.34387383
+ pdiblc2 = 0.0089064378
+ pdiblcb = -0.035822256
+ drout = 0.47767008
+ pscbe1 = 7.9223209e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_23}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_23}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.24044135+sky130_fd_pr__nfet_01v8__kt1_diff_23}
+ kt2 = -0.029182241
+ at = 58808.073
+ ute = 0.0
+ ua1 = 1.8137456e-9
+ ub1 = -6.1118594e-19
+ uc1 = 1.4013253e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.24 nmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.48265+sky130_fd_pr__nfet_01v8__vth0_diff_24+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.88719062
+ k2 = {-0.12944+sky130_fd_pr__nfet_01v8__k2_diff_24}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {136940+sky130_fd_pr__nfet_01v8__vsat_diff_24}
+ ua = {-7.6981e-010+sky130_fd_pr__nfet_01v8__ua_diff_24}
+ ub = {1.8891e-018+sky130_fd_pr__nfet_01v8__ub_diff_24}
+ uc = 8.1344e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_24}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.035567+sky130_fd_pr__nfet_01v8__u0_diff_24}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_24}
+ keta = {-0.044024+sky130_fd_pr__nfet_01v8__keta_diff_24}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_24}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_24}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_24}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.14634+sky130_fd_pr__nfet_01v8__voff_diff_24+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.7368+sky130_fd_pr__nfet_01v8__nfactor_diff_24+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_24}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.037587994+sky130_fd_pr__nfet_01v8__eta0_diff_24}
+ etab = -0.025196
+ dsub = 0.39524783
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.3933+sky130_fd_pr__nfet_01v8__pclm_diff_24}
+ pdiblc1 = 0.37540586
+ pdiblc2 = 0.0092926225
+ pdiblcb = -0.10619144
+ drout = 0.80296042
+ pscbe1 = 7.9758201e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7248e-6
+ alpha1 = 0.67137
+ beta0 = 18.392
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_24}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_24}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27282685+sky130_fd_pr__nfet_01v8__kt1_diff_24}
+ kt2 = -0.035936577
+ at = 44113.722
+ ute = -1.8337678
+ ua1 = -5.4118864e-10
+ ub1 = 7.8192473e-19
+ uc1 = 9.8973497e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.25 nmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.53379+sky130_fd_pr__nfet_01v8__vth0_diff_25+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.7651852
+ k2 = {-0.093246775+sky130_fd_pr__nfet_01v8__k2_diff_25}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {138200+sky130_fd_pr__nfet_01v8__vsat_diff_25}
+ ua = {-2.1195046e-009+sky130_fd_pr__nfet_01v8__ua_diff_25}
+ ub = {2.388e-018+sky130_fd_pr__nfet_01v8__ub_diff_25}
+ uc = 4.7656998e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_25}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.018279679+sky130_fd_pr__nfet_01v8__u0_diff_25}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_25}
+ keta = {-0.03233914+sky130_fd_pr__nfet_01v8__keta_diff_25}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.01953125+sky130_fd_pr__nfet_01v8__ags_diff_25}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_25}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_25}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.14315115+sky130_fd_pr__nfet_01v8__voff_diff_25+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.7329074+sky130_fd_pr__nfet_01v8__nfactor_diff_25+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_25}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.49+sky130_fd_pr__nfet_01v8__eta0_diff_25}
+ etab = -0.0010980414
+ dsub = 0.53787594
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.42537+sky130_fd_pr__nfet_01v8__pclm_diff_25}
+ pdiblc1 = 0.49955094
+ pdiblc2 = 0.0025320601
+ pdiblcb = -0.025
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.5e-6
+ alpha1 = 0.85
+ beta0 = 19.404
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_25}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_25}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27356256+sky130_fd_pr__nfet_01v8__kt1_diff_25}
+ kt2 = -0.026436448
+ at = 27185.354
+ ute = -0.64193177
+ ua1 = 1.6863756e-9
+ ub1 = -8.6491606e-19
+ uc1 = 7.9489697e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.26 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.58492159+sky130_fd_pr__nfet_01v8__vth0_diff_26+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47758412
+ k2 = {-0.0092134864+sky130_fd_pr__nfet_01v8__k2_diff_26}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {124450+sky130_fd_pr__nfet_01v8__vsat_diff_26}
+ ua = {-1.5528769e-009+sky130_fd_pr__nfet_01v8__ua_diff_26}
+ ub = {2.1949e-018+sky130_fd_pr__nfet_01v8__ub_diff_26}
+ uc = 8.1535e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_26}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.024442+sky130_fd_pr__nfet_01v8__u0_diff_26}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_26}
+ keta = {-0.021959431+sky130_fd_pr__nfet_01v8__keta_diff_26}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_26}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_26}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_26}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.13972753+sky130_fd_pr__nfet_01v8__voff_diff_26+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.5922074+sky130_fd_pr__nfet_01v8__nfactor_diff_26+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_26}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.49+sky130_fd_pr__nfet_01v8__eta0_diff_26}
+ etab = -0.0003125
+ dsub = 0.3565784
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.42387+sky130_fd_pr__nfet_01v8__pclm_diff_26}
+ pdiblc1 = 0.87848679
+ pdiblc2 = 0.0030018173
+ pdiblcb = -0.025
+ drout = 0.91727235
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_26}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_26}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27851007+sky130_fd_pr__nfet_01v8__kt1_diff_26}
+ kt2 = -0.036334685
+ at = 53841.958
+ ute = -1.4717587
+ ua1 = 1.0329816e-9
+ ub1 = -1.136817e-18
+ uc1 = -1.275902e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.27 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.56984+sky130_fd_pr__nfet_01v8__vth0_diff_27+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.58363587
+ k2 = {-0.050449684+sky130_fd_pr__nfet_01v8__k2_diff_27}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {100300+sky130_fd_pr__nfet_01v8__vsat_diff_27}
+ ua = {-1.448307e-009+sky130_fd_pr__nfet_01v8__ua_diff_27}
+ ub = {2.2568e-018+sky130_fd_pr__nfet_01v8__ub_diff_27}
+ uc = 6.0873e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_27}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.027403+sky130_fd_pr__nfet_01v8__u0_diff_27}
+ a0 = {1.02+sky130_fd_pr__nfet_01v8__a0_diff_27}
+ keta = {-0.065071813+sky130_fd_pr__nfet_01v8__keta_diff_27}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.95+sky130_fd_pr__nfet_01v8__ags_diff_27}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_27}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_27}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.12063615+sky130_fd_pr__nfet_01v8__voff_diff_27+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.6637647+sky130_fd_pr__nfet_01v8__nfactor_diff_27+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_27}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.00253125+sky130_fd_pr__nfet_01v8__eta0_diff_27}
+ etab = -0.0003125
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.39168+sky130_fd_pr__nfet_01v8__pclm_diff_27}
+ pdiblc1 = 0.7071625
+ pdiblc2 = 0.004011417
+ pdiblcb = -0.00019159217
+ drout = 0.26
+ pscbe1 = 2.6107456e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.64e-6
+ alpha1 = 0.884
+ beta0 = 16.632
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_27}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_27}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27269+sky130_fd_pr__nfet_01v8__kt1_diff_27}
+ kt2 = -0.026386792
+ at = 63366.0
+ ute = -0.88681922
+ ua1 = 2.2042059e-9
+ ub1 = -1.4677553e-18
+ uc1 = 5.5867248e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.28 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.53889+sky130_fd_pr__nfet_01v8__vth0_diff_28+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.5498852
+ k2 = {-0.038377686+sky130_fd_pr__nfet_01v8__k2_diff_28}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_28}
+ ua = {-9.3056317e-010+sky130_fd_pr__nfet_01v8__ua_diff_28}
+ ub = {1.8431e-018+sky130_fd_pr__nfet_01v8__ub_diff_28}
+ uc = 7.4314e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_28}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.031624+sky130_fd_pr__nfet_01v8__u0_diff_28}
+ a0 = {1.1868+sky130_fd_pr__nfet_01v8__a0_diff_28}
+ keta = {-0.00012732+sky130_fd_pr__nfet_01v8__keta_diff_28}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.60805+sky130_fd_pr__nfet_01v8__ags_diff_28}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_28}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_28}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.10191764+sky130_fd_pr__nfet_01v8__voff_diff_28+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_28+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_28}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.0005+sky130_fd_pr__nfet_01v8__eta0_diff_28}
+ etab = -0.00050069107
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.55915+sky130_fd_pr__nfet_01v8__pclm_diff_28}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0048124934
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_28}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_28}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.32398+sky130_fd_pr__nfet_01v8__kt1_diff_28}
+ kt2 = -0.046448585
+ at = 114940.0
+ ute = -1.7149
+ ua1 = 4.8534e-10
+ ub1 = -5.6531e-19
+ uc1 = 3.6436037e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.29 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.53475+sky130_fd_pr__nfet_01v8__vth0_diff_29+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 0.55001325
+ k2 = {-0.035329605+sky130_fd_pr__nfet_01v8__k2_diff_29}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_29}
+ ua = {-7.5728632e-010+sky130_fd_pr__nfet_01v8__ua_diff_29}
+ ub = {1.6878e-018+sky130_fd_pr__nfet_01v8__ub_diff_29}
+ uc = 4.2895e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_29}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.033+sky130_fd_pr__nfet_01v8__u0_diff_29}
+ a0 = {1.26+sky130_fd_pr__nfet_01v8__a0_diff_29}
+ keta = {-0.0019819+sky130_fd_pr__nfet_01v8__keta_diff_29}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.39508+sky130_fd_pr__nfet_01v8__ags_diff_29}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_29}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_29}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.10164906+sky130_fd_pr__nfet_01v8__voff_diff_29+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_29+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_29}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_29}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.58702+sky130_fd_pr__nfet_01v8__pclm_diff_29}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.003090586
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_29}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_29}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.31514+sky130_fd_pr__nfet_01v8__kt1_diff_29}
+ kt2 = -0.046434757
+ at = 140000.0
+ ute = -1.8532
+ ua1 = 1.7906e-10
+ ub1 = -3.8177e-19
+ uc1 = 3.0357419e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.30 nmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.5214+sky130_fd_pr__nfet_01v8__vth0_diff_30+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.54086565
+ k2 = {-0.031031091+sky130_fd_pr__nfet_01v8__k2_diff_30}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_30}
+ ua = {-7.6156997e-010+sky130_fd_pr__nfet_01v8__ua_diff_30}
+ ub = {1.7377e-018+sky130_fd_pr__nfet_01v8__ub_diff_30}
+ uc = 4.9242e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_30}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.033074+sky130_fd_pr__nfet_01v8__u0_diff_30}
+ a0 = {1.32+sky130_fd_pr__nfet_01v8__a0_diff_30}
+ keta = {-0.0087946+sky130_fd_pr__nfet_01v8__keta_diff_30}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.40535+sky130_fd_pr__nfet_01v8__ags_diff_30}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_30}
+ b1 = {2.1073424e-024+sky130_fd_pr__nfet_01v8__b1_diff_30}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.1052686+sky130_fd_pr__nfet_01v8__voff_diff_30+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_30+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_30}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_30}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.026316+sky130_fd_pr__nfet_01v8__pclm_diff_30}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0030734587
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.5467416e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_30}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_30}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.31303+sky130_fd_pr__nfet_01v8__kt1_diff_30}
+ kt2 = -0.045313337
+ at = 140000.0
+ ute = -1.8134
+ ua1 = 3.7602e-10
+ ub1 = -6.3962e-19
+ uc1 = 1.5829713e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.31 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.43529+sky130_fd_pr__nfet_01v8__vth0_diff_31+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 0.90272985
+ k2 = {-0.12855+sky130_fd_pr__nfet_01v8__k2_diff_31}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {159360+sky130_fd_pr__nfet_01v8__vsat_diff_31}
+ ua = {-2.3936e-009+sky130_fd_pr__nfet_01v8__ua_diff_31}
+ ub = {2.7296e-018+sky130_fd_pr__nfet_01v8__ub_diff_31}
+ uc = 5.3128e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_31}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.015121+sky130_fd_pr__nfet_01v8__u0_diff_31}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_31}
+ keta = {0.022506+sky130_fd_pr__nfet_01v8__keta_diff_31}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_31}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_31}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_31}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.21786+sky130_fd_pr__nfet_01v8__voff_diff_31+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.9783+sky130_fd_pr__nfet_01v8__nfactor_diff_31+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_31}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.0007818+sky130_fd_pr__nfet_01v8__eta0_diff_31}
+ etab = -0.042588
+ dsub = 0.32653
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.16949+sky130_fd_pr__nfet_01v8__pclm_diff_31}
+ pdiblc1 = 0.38670965
+ pdiblc2 = 0.0095519
+ pdiblcb = -9.5889633e-6
+ drout = 0.53658367
+ pscbe1 = 7.9053558e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_31}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_31}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.21542+sky130_fd_pr__nfet_01v8__kt1_diff_31}
+ kt2 = -0.029433449
+ at = 32729.0
+ ute = 0.0
+ ua1 = 1.986e-9
+ ub1 = -5.3915e-19
+ uc1 = 1.5881061e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.32 nmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.48847+sky130_fd_pr__nfet_01v8__vth0_diff_32+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.88672771
+ k2 = {-0.13044547+sky130_fd_pr__nfet_01v8__k2_diff_32}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {148510+sky130_fd_pr__nfet_01v8__vsat_diff_32}
+ ua = {-7.8712e-010+sky130_fd_pr__nfet_01v8__ua_diff_32}
+ ub = {1.9242e-018+sky130_fd_pr__nfet_01v8__ub_diff_32}
+ uc = 8.6399e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_32}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.035452+sky130_fd_pr__nfet_01v8__u0_diff_32}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_32}
+ keta = {-0.039244+sky130_fd_pr__nfet_01v8__keta_diff_32}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_32}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_32}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_32}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.15486+sky130_fd_pr__nfet_01v8__voff_diff_32+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.6549+sky130_fd_pr__nfet_01v8__nfactor_diff_32+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_32}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.030982769+sky130_fd_pr__nfet_01v8__eta0_diff_32}
+ etab = -0.028357517
+ dsub = 0.3989415
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.28643+sky130_fd_pr__nfet_01v8__pclm_diff_32}
+ pdiblc1 = 0.37487423
+ pdiblc2 = 0.0088295033
+ pdiblcb = -0.086356118
+ drout = 0.71690147
+ pscbe1 = 7.9589649e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.802e-9
+ alpha1 = 1.1911
+ beta0 = 15.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_32}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_32}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25912854+sky130_fd_pr__nfet_01v8__kt1_diff_32}
+ kt2 = -0.036161033
+ at = 35966.431
+ ute = -1.8244516
+ ua1 = -5.5496972e-10
+ ub1 = 9.1703372e-19
+ uc1 = 1.3163208e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.33 nmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.53303+sky130_fd_pr__nfet_01v8__vth0_diff_33+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.76175334
+ k2 = {-0.092823426+sky130_fd_pr__nfet_01v8__k2_diff_33}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {141560+sky130_fd_pr__nfet_01v8__vsat_diff_33}
+ ua = {-2.1372071e-009+sky130_fd_pr__nfet_01v8__ua_diff_33}
+ ub = {2.5013e-018+sky130_fd_pr__nfet_01v8__ub_diff_33}
+ uc = 8.4588e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_33}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.018858+sky130_fd_pr__nfet_01v8__u0_diff_33}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_33}
+ keta = {-0.038557533+sky130_fd_pr__nfet_01v8__keta_diff_33}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.019531+sky130_fd_pr__nfet_01v8__ags_diff_33}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_33}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_33}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.1423314+sky130_fd_pr__nfet_01v8__voff_diff_33+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8066026+sky130_fd_pr__nfet_01v8__nfactor_diff_33+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_33}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.49+sky130_fd_pr__nfet_01v8__eta0_diff_33}
+ etab = -0.00088983339
+ dsub = 0.55793099
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.41199+sky130_fd_pr__nfet_01v8__pclm_diff_33}
+ pdiblc1 = 0.11815701
+ pdiblc2 = 0.002539823
+ pdiblcb = -0.225
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.64e-6
+ alpha1 = 0.85
+ beta0 = 19.127
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_33}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_33}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.29166204+sky130_fd_pr__nfet_01v8__kt1_diff_33}
+ kt2 = -0.039951188
+ at = 25924.417
+ ute = -0.86888901
+ ua1 = 1.4604853e-9
+ ub1 = -7.67306e-19
+ uc1 = 9.0064279e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.34 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.58177+sky130_fd_pr__nfet_01v8__vth0_diff_34+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.48574418
+ k2 = {-0.010465693+sky130_fd_pr__nfet_01v8__k2_diff_34}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {115210+sky130_fd_pr__nfet_01v8__vsat_diff_34}
+ ua = {-1.6072627e-009+sky130_fd_pr__nfet_01v8__ua_diff_34}
+ ub = {2.2467e-018+sky130_fd_pr__nfet_01v8__ub_diff_34}
+ uc = 8.2749e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_34}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.024026+sky130_fd_pr__nfet_01v8__u0_diff_34}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_34}
+ keta = {-0.026851+sky130_fd_pr__nfet_01v8__keta_diff_34}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_34}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_34}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_34}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.13427734+sky130_fd_pr__nfet_01v8__voff_diff_34+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.7157106+sky130_fd_pr__nfet_01v8__nfactor_diff_34+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_34}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.49+sky130_fd_pr__nfet_01v8__eta0_diff_34}
+ etab = -0.0003125
+ dsub = 0.39550151
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.5366+sky130_fd_pr__nfet_01v8__pclm_diff_34}
+ pdiblc1 = 1.0
+ pdiblc2 = 0.0034253023
+ pdiblcb = -0.025
+ drout = 0.49875239
+ pscbe1 = 5.6082016e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.0e-6
+ alpha1 = 0.85
+ beta0 = 18.8
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_34}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_34}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27675+sky130_fd_pr__nfet_01v8__kt1_diff_34}
+ kt2 = -0.036077934
+ at = 53428.0
+ ute = -1.4271
+ ua1 = 1.1226477e-9
+ ub1 = -1.1992841e-18
+ uc1 = -1.3721851e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.35 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.53913942+sky130_fd_pr__nfet_01v8__vth0_diff_35+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.58562329
+ k2 = {-0.056895912+sky130_fd_pr__nfet_01v8__k2_diff_35}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {176000+sky130_fd_pr__nfet_01v8__vsat_diff_35}
+ ua = {-1.2391262e-009+sky130_fd_pr__nfet_01v8__ua_diff_35}
+ ub = {1.8409e-018+sky130_fd_pr__nfet_01v8__ub_diff_35}
+ uc = 4.2541e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_35}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.028539+sky130_fd_pr__nfet_01v8__u0_diff_35}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_35}
+ keta = {0.017793861+sky130_fd_pr__nfet_01v8__keta_diff_35}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.20227+sky130_fd_pr__nfet_01v8__ags_diff_35}
+ b0 = {-8.9909e-008+sky130_fd_pr__nfet_01v8__b0_diff_35}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_35}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.11956669+sky130_fd_pr__nfet_01v8__voff_diff_35+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.5286687+sky130_fd_pr__nfet_01v8__nfactor_diff_35+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_35}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.00253125+sky130_fd_pr__nfet_01v8__eta0_diff_35}
+ etab = -0.0003125
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {1.0354+sky130_fd_pr__nfet_01v8__pclm_diff_35}
+ pdiblc1 = 0.58940551
+ pdiblc2 = 0.0058383177
+ pdiblcb = -0.025
+ drout = 0.65422372
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_35}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_35}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.29597636+sky130_fd_pr__nfet_01v8__kt1_diff_35}
+ kt2 = -0.02645877
+ at = 130000.0
+ ute = -0.71912805
+ ua1 = 2.1943519e-9
+ ub1 = -1.3628408e-18
+ uc1 = 4.7561934e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.36 nmos
* DC IV MOS Parameters
+ lmin = 1.9995e-05 lmax = 2.0005e-05 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.49711+sky130_fd_pr__nfet_01v8__vth0_diff_36+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = {-0.041590846+sky130_fd_pr__nfet_01v8__k2_diff_36}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_36}
+ ua = {-1.0612493e-009+sky130_fd_pr__nfet_01v8__ua_diff_36}
+ ub = {1.7139e-018+sky130_fd_pr__nfet_01v8__ub_diff_36}
+ uc = 4.8537e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_36}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.027964+sky130_fd_pr__nfet_01v8__u0_diff_36}
+ a0 = {1.3626+sky130_fd_pr__nfet_01v8__a0_diff_36}
+ keta = {-0.0045466+sky130_fd_pr__nfet_01v8__keta_diff_36}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.34488+sky130_fd_pr__nfet_01v8__ags_diff_36}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_36}
+ b1 = {2.1073424e-024+sky130_fd_pr__nfet_01v8__b1_diff_36}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_diff_36+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_36+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_36}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_36}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.016875+sky130_fd_pr__nfet_01v8__pclm_diff_36}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.25e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_36}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_36}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.28638+sky130_fd_pr__nfet_01v8__kt1_diff_36}
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.37 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.55051256+sky130_fd_pr__nfet_01v8__vth0_diff_37+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.6038851
+ k2 = {-0.063708056+sky130_fd_pr__nfet_01v8__k2_diff_37}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {148000+sky130_fd_pr__nfet_01v8__vsat_diff_37}
+ ua = {-7.4248288e-010+sky130_fd_pr__nfet_01v8__ua_diff_37}
+ ub = {1.5791e-018+sky130_fd_pr__nfet_01v8__ub_diff_37}
+ uc = 4.5455e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_37}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.033776+sky130_fd_pr__nfet_01v8__u0_diff_37}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_37}
+ keta = {0.017925112+sky130_fd_pr__nfet_01v8__keta_diff_37}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.26838+sky130_fd_pr__nfet_01v8__ags_diff_37}
+ b0 = {-6e-008+sky130_fd_pr__nfet_01v8__b0_diff_37}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_37}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.10864023+sky130_fd_pr__nfet_01v8__voff_diff_37+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_37+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_37}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_37}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {1.7974+sky130_fd_pr__nfet_01v8__pclm_diff_37}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.01341528
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_37}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_37}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.32201+sky130_fd_pr__nfet_01v8__kt1_diff_37}
+ kt2 = -0.030441716
+ at = 140000.0
+ ute = -1.1848
+ ua1 = 1.4932e-9
+ ub1 = -8.92e-19
+ uc1 = 4.5225072e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.38 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.53566+sky130_fd_pr__nfet_01v8__vth0_diff_38+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 0.56269175
+ k2 = {-0.049175583+sky130_fd_pr__nfet_01v8__k2_diff_38}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_38}
+ ua = {-6.1895011e-010+sky130_fd_pr__nfet_01v8__ua_diff_38}
+ ub = {1.3523e-018+sky130_fd_pr__nfet_01v8__ub_diff_38}
+ uc = 2.0e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_38}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.032099+sky130_fd_pr__nfet_01v8__u0_diff_38}
+ a0 = {1.17+sky130_fd_pr__nfet_01v8__a0_diff_38}
+ keta = {0.0024561+sky130_fd_pr__nfet_01v8__keta_diff_38}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.35354+sky130_fd_pr__nfet_01v8__ags_diff_38}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_38}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_38}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.1101223+sky130_fd_pr__nfet_01v8__voff_diff_38+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_38+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_38}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_38}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.51494+sky130_fd_pr__nfet_01v8__pclm_diff_38}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0063461484
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_38}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_38}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.3138+sky130_fd_pr__nfet_01v8__kt1_diff_38}
+ kt2 = -0.043698517
+ at = 140000.0
+ ute = -1.4002
+ ua1 = 5.7852e-10
+ ub1 = -4.1255e-19
+ uc1 = 5.1716116e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.39 nmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.51412+sky130_fd_pr__nfet_01v8__vth0_diff_39+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.585057
+ k2 = {-0.049134061+sky130_fd_pr__nfet_01v8__k2_diff_39}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_39}
+ ua = {-9.2975583e-010+sky130_fd_pr__nfet_01v8__ua_diff_39}
+ ub = {1.6982e-018+sky130_fd_pr__nfet_01v8__ub_diff_39}
+ uc = 2.6301e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_39}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.029912+sky130_fd_pr__nfet_01v8__u0_diff_39}
+ a0 = {1.188+sky130_fd_pr__nfet_01v8__a0_diff_39}
+ keta = {-0.0084252+sky130_fd_pr__nfet_01v8__keta_diff_39}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.38014+sky130_fd_pr__nfet_01v8__ags_diff_39}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_39}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_39}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.11808229+sky130_fd_pr__nfet_01v8__voff_diff_39+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_39+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_39}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_39}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.083531+sky130_fd_pr__nfet_01v8__pclm_diff_39}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0026381856
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.6297212e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_39}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_39}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.29822+sky130_fd_pr__nfet_01v8__kt1_diff_39}
+ kt2 = -0.031096922
+ at = 155000.0
+ ute = -1.1026
+ ua1 = 1.4885e-9
+ ub1 = -1.0524e-18
+ uc1 = 1.9763869e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.40 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.42664+sky130_fd_pr__nfet_01v8__vth0_diff_40+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.14006+sky130_fd_pr__nfet_01v8__k2_diff_40}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {193330+sky130_fd_pr__nfet_01v8__vsat_diff_40}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_40}
+ ub = {2.0811e-018+sky130_fd_pr__nfet_01v8__ub_diff_40}
+ uc = 6.8253e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_40}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.029497+sky130_fd_pr__nfet_01v8__u0_diff_40}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_40}
+ keta = {-0.0924+sky130_fd_pr__nfet_01v8__keta_diff_40}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_40}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_40}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_40}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_40+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.612+sky130_fd_pr__nfet_01v8__nfactor_diff_40+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_40}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0+sky130_fd_pr__nfet_01v8__eta0_diff_40}
+ etab = -0.043998
+ dsub = 0.62373
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.14377+sky130_fd_pr__nfet_01v8__pclm_diff_40}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.85
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_40}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_40}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.24096074+sky130_fd_pr__nfet_01v8__kt1_diff_40}
+ kt2 = -0.028878939
+ at = 53720.487
+ ute = -1.2190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.41 nmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.48404+sky130_fd_pr__nfet_01v8__vth0_diff_41+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.14006+sky130_fd_pr__nfet_01v8__k2_diff_41}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {198330+sky130_fd_pr__nfet_01v8__vsat_diff_41}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_41}
+ ub = {2.1643e-018+sky130_fd_pr__nfet_01v8__ub_diff_41}
+ uc = 9.1459e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_41}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.031005+sky130_fd_pr__nfet_01v8__u0_diff_41}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_41}
+ keta = {-0.068376+sky130_fd_pr__nfet_01v8__keta_diff_41}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_41}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_41}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_41}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_41+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {0.87048+sky130_fd_pr__nfet_01v8__nfactor_diff_41+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_41}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0+sky130_fd_pr__nfet_01v8__eta0_diff_41}
+ etab = -0.043998
+ dsub = 0.62373
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.18115+sky130_fd_pr__nfet_01v8__pclm_diff_41}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.16e-8
+ alpha1 = 0.85
+ beta0 = 14.4
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_41}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_41}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.22096074+sky130_fd_pr__nfet_01v8__kt1_diff_41}
+ kt2 = -0.028878939
+ at = 43720.487
+ ute = -1.2790432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.42 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.55302+sky130_fd_pr__nfet_01v8__vth0_diff_42+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57549796
+ k2 = {-0.056325504+sky130_fd_pr__nfet_01v8__k2_diff_42}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {193940+sky130_fd_pr__nfet_01v8__vsat_diff_42}
+ ua = {-1.1764338e-009+sky130_fd_pr__nfet_01v8__ua_diff_42}
+ ub = {1.706e-018+sky130_fd_pr__nfet_01v8__ub_diff_42}
+ uc = 4.4038254e-12
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_42}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.02858942+sky130_fd_pr__nfet_01v8__u0_diff_42}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_42}
+ keta = {-0.0017502917+sky130_fd_pr__nfet_01v8__keta_diff_42}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.01953125+sky130_fd_pr__nfet_01v8__ags_diff_42}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_42}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_42}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.1331126+sky130_fd_pr__nfet_01v8__voff_diff_42+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.7358334+sky130_fd_pr__nfet_01v8__nfactor_diff_42+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_42}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.49+sky130_fd_pr__nfet_01v8__eta0_diff_42}
+ etab = -0.0003125
+ dsub = 0.30522325
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62116627+sky130_fd_pr__nfet_01v8__pclm_diff_42}
+ pdiblc1 = 0.49968287
+ pdiblc2 = 0.0013250286
+ pdiblcb = -0.025
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.0e-7
+ alpha1 = 0.85
+ beta0 = 15.6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_42}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_42}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.30582115+sky130_fd_pr__nfet_01v8__kt1_diff_42}
+ kt2 = -0.049881868
+ at = 0.0
+ ute = -1.4845028
+ ua1 = 3.7866659e-10
+ ub1 = 5.2996898e-20
+ uc1 = 1.0632025e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.43 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.54988+sky130_fd_pr__nfet_01v8__vth0_diff_43+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55418882
+ k2 = {-0.045978853+sky130_fd_pr__nfet_01v8__k2_diff_43}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {83416+sky130_fd_pr__nfet_01v8__vsat_diff_43}
+ ua = {-1.1390319e-009+sky130_fd_pr__nfet_01v8__ua_diff_43}
+ ub = {1.742e-018+sky130_fd_pr__nfet_01v8__ub_diff_43}
+ uc = 3.9553e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_43}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.02797+sky130_fd_pr__nfet_01v8__u0_diff_43}
+ a0 = {1.2+sky130_fd_pr__nfet_01v8__a0_diff_43}
+ keta = {-0.062678008+sky130_fd_pr__nfet_01v8__keta_diff_43}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_43}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_43}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_43}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.1346663+sky130_fd_pr__nfet_01v8__voff_diff_43+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.3985224+sky130_fd_pr__nfet_01v8__nfactor_diff_43+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_43}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.00253125+sky130_fd_pr__nfet_01v8__eta0_diff_43}
+ etab = -0.084375
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.87034+sky130_fd_pr__nfet_01v8__pclm_diff_43}
+ pdiblc1 = 0.35436836
+ pdiblc2 = 0.0046946379
+ pdiblcb = -0.00019150181
+ drout = 0.91970352
+ pscbe1 = 7.3389715e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.52e-6
+ alpha1 = 0.85
+ beta0 = 17.464
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_43}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_43}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27465702+sky130_fd_pr__nfet_01v8__kt1_diff_43}
+ kt2 = -0.027125854
+ at = 62688.03
+ ute = -1.0746097
+ ua1 = 1.2815636e-9
+ ub1 = -6.7036132e-19
+ uc1 = 4.1015542e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.44 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.54039+sky130_fd_pr__nfet_01v8__vth0_diff_44+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57309884
+ k2 = {-0.05049203+sky130_fd_pr__nfet_01v8__k2_diff_44}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_44}
+ ua = {-4.4055851e-010+sky130_fd_pr__nfet_01v8__ua_diff_44}
+ ub = {1.4e-018+sky130_fd_pr__nfet_01v8__ub_diff_44}
+ uc = 5.079e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_44}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.035815+sky130_fd_pr__nfet_01v8__u0_diff_44}
+ a0 = {0.8448+sky130_fd_pr__nfet_01v8__a0_diff_44}
+ keta = {0.0050203+sky130_fd_pr__nfet_01v8__keta_diff_44}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.47645+sky130_fd_pr__nfet_01v8__ags_diff_44}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_44}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_44}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.09931841+sky130_fd_pr__nfet_01v8__voff_diff_44+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_44+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_44}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.0005+sky130_fd_pr__nfet_01v8__eta0_diff_44}
+ etab = -0.0005
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.50564+sky130_fd_pr__nfet_01v8__pclm_diff_44}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0071800746
+ pdiblcb = -0.0125
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_44}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_44}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.33382+sky130_fd_pr__nfet_01v8__kt1_diff_44}
+ kt2 = -0.048264621
+ at = 109370.0
+ ute = -1.7304
+ ua1 = -1.5662e-10
+ ub1 = 1.5093e-19
+ uc1 = 5.6582773e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.45 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.5364+sky130_fd_pr__nfet_01v8__vth0_diff_45+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56608288
+ k2 = {-0.045363238+sky130_fd_pr__nfet_01v8__k2_diff_45}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_45}
+ ua = {-5.7533961e-010+sky130_fd_pr__nfet_01v8__ua_diff_45}
+ ub = {1.4937e-018+sky130_fd_pr__nfet_01v8__ub_diff_45}
+ uc = 4.3137e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_45}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.033505+sky130_fd_pr__nfet_01v8__u0_diff_45}
+ a0 = {1.23+sky130_fd_pr__nfet_01v8__a0_diff_45}
+ keta = {0.0027556+sky130_fd_pr__nfet_01v8__keta_diff_45}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.40117+sky130_fd_pr__nfet_01v8__ags_diff_45}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_45}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_45}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.11839262+sky130_fd_pr__nfet_01v8__voff_diff_45+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.7745196+sky130_fd_pr__nfet_01v8__nfactor_diff_45+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_45}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_45}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.81282+sky130_fd_pr__nfet_01v8__pclm_diff_45}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0048130092
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.1120295e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_45}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_45}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.29604+sky130_fd_pr__nfet_01v8__kt1_diff_45}
+ kt2 = -0.031412161
+ at = 140000.0
+ ute = -1.2994
+ ua1 = 9.9875e-10
+ ub1 = -6.725e-19
+ uc1 = 3.2355466e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.46 nmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.52187+sky130_fd_pr__nfet_01v8__vth0_diff_46+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.50132234
+ k2 = {-0.017423723+sky130_fd_pr__nfet_01v8__k2_diff_46}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80000+sky130_fd_pr__nfet_01v8__vsat_diff_46}
+ ua = {-7.7745124e-010+sky130_fd_pr__nfet_01v8__ua_diff_46}
+ ub = {1.4645e-018+sky130_fd_pr__nfet_01v8__ub_diff_46}
+ uc = 2.6318e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_46}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.030087+sky130_fd_pr__nfet_01v8__u0_diff_46}
+ a0 = {1.32+sky130_fd_pr__nfet_01v8__a0_diff_46}
+ keta = {-0.0073844+sky130_fd_pr__nfet_01v8__keta_diff_46}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.38101+sky130_fd_pr__nfet_01v8__ags_diff_46}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_46}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_46}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.11819485+sky130_fd_pr__nfet_01v8__voff_diff_46+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.8+sky130_fd_pr__nfet_01v8__nfactor_diff_46+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_46}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8__eta0_diff_46}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.056875+sky130_fd_pr__nfet_01v8__pclm_diff_46}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0015751675
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.7499921e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_46}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_46}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.29114+sky130_fd_pr__nfet_01v8__kt1_diff_46}
+ kt2 = -0.020571319
+ at = 140000.0
+ ute = -1.2651
+ ua1 = 1.2581e-9
+ ub1 = -8.5051e-19
+ uc1 = -1.9578625e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.47 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.46461+sky130_fd_pr__nfet_01v8__vth0_diff_47+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.13467+sky130_fd_pr__nfet_01v8__k2_diff_47}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {185700+sky130_fd_pr__nfet_01v8__vsat_diff_47}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_47}
+ ub = {2.3194e-018+sky130_fd_pr__nfet_01v8__ub_diff_47}
+ uc = 8.7504e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_47}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.029597+sky130_fd_pr__nfet_01v8__u0_diff_47}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_47}
+ keta = {-0.027+sky130_fd_pr__nfet_01v8__keta_diff_47}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_47}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_47}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_47}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_47+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {2.015+sky130_fd_pr__nfet_01v8__nfactor_diff_47+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_47}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0.00069413878+sky130_fd_pr__nfet_01v8__eta0_diff_47}
+ etab = -0.043998
+ dsub = 0.45862506
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.16337+sky130_fd_pr__nfet_01v8__pclm_diff_47}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.85
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_47}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_47}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.24096074+sky130_fd_pr__nfet_01v8__kt1_diff_47}
+ kt2 = -0.028878939
+ at = 53720.487
+ ute = -1.2550432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.48 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.57828+sky130_fd_pr__nfet_01v8__vth0_diff_48+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47498405
+ k2 = {-0.011809992+sky130_fd_pr__nfet_01v8__k2_diff_48}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {184270+sky130_fd_pr__nfet_01v8__vsat_diff_48}
+ ua = {-1.4557395e-009+sky130_fd_pr__nfet_01v8__ua_diff_48}
+ ub = {1.9002e-018+sky130_fd_pr__nfet_01v8__ub_diff_48}
+ uc = 5.2537e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_48}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.023543+sky130_fd_pr__nfet_01v8__u0_diff_48}
+ a0 = {1.3846+sky130_fd_pr__nfet_01v8__a0_diff_48}
+ keta = {-0.0071133131+sky130_fd_pr__nfet_01v8__keta_diff_48}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {0.15625+sky130_fd_pr__nfet_01v8__ags_diff_48}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_48}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_48}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.14363643+sky130_fd_pr__nfet_01v8__voff_diff_48+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {1.3263601+sky130_fd_pr__nfet_01v8__nfactor_diff_48+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_48}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ eta0 = {0.49+sky130_fd_pr__nfet_01v8__eta0_diff_48}
+ etab = -0.000625
+ dsub = 0.31030713
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.45181+sky130_fd_pr__nfet_01v8__pclm_diff_48}
+ pdiblc1 = 0.033031793
+ pdiblc2 = 4.6437666e-5
+ pdiblcb = -0.09460521
+ drout = 0.9999999
+ pscbe1 = 4.3694701e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.9e-6
+ alpha1 = 0.85
+ beta0 = 18.018
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_48}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_48}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27894958+sky130_fd_pr__nfet_01v8__kt1_diff_48}
+ kt2 = -0.0367186
+ at = 10655.26
+ ute = -1.3102789
+ ua1 = 8.3166957e-10
+ ub1 = -6.31879e-19
+ uc1 = 5.7404281e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.49 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 6.35e-07 wmax = 6.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.45263+sky130_fd_pr__nfet_01v8__vth0_diff_49+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.13467+sky130_fd_pr__nfet_01v8__k2_diff_49}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {170440+sky130_fd_pr__nfet_01v8__vsat_diff_49}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_49}
+ ub = {2.1338e-018+sky130_fd_pr__nfet_01v8__ub_diff_49}
+ uc = 7.7004e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_49}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.030197+sky130_fd_pr__nfet_01v8__u0_diff_49}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_49}
+ keta = {-0.027+sky130_fd_pr__nfet_01v8__keta_diff_49}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_49}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_49}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_49}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_49+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {2.015+sky130_fd_pr__nfet_01v8__nfactor_diff_49+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_49}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0+sky130_fd_pr__nfet_01v8__eta0_diff_49}
+ etab = -0.043998
+ dsub = 0.45863
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.18297+sky130_fd_pr__nfet_01v8__pclm_diff_49}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.85
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_49}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_49}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.23096074+sky130_fd_pr__nfet_01v8__kt1_diff_49}
+ kt2 = -0.028878939
+ at = 53720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.50 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 8.35e-07 wmax = 8.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.1932e-008+sky130_fd_pr__nfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1859e-008+sky130_fd_pr__nfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -1.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8__rshn_mult}
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.48208+sky130_fd_pr__nfet_01v8__vth0_diff_50+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.12659+sky130_fd_pr__nfet_01v8__k2_diff_50}
+ k3 = 2.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ w0 = 0.0
+ k3b = 0.54
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {179460+sky130_fd_pr__nfet_01v8__vsat_diff_50}
+ ua = {-1.1926e-009+sky130_fd_pr__nfet_01v8__ua_diff_50}
+ ub = {2.1338e-018+sky130_fd_pr__nfet_01v8__ub_diff_50}
+ uc = 7.7004e-11
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_50}
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
+ u0 = {0.029027+sky130_fd_pr__nfet_01v8__u0_diff_50}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_50}
+ keta = {-0.027+sky130_fd_pr__nfet_01v8__keta_diff_50}
+ a1 = 0.0
+ a2 = 0.42385546
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_50}
+ b0 = {0+sky130_fd_pr__nfet_01v8__b0_diff_50}
+ b1 = {0+sky130_fd_pr__nfet_01v8__b1_diff_50}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_50+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {2.015+sky130_fd_pr__nfet_01v8__nfactor_diff_50+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8__tvoff_diff_50}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ eta0 = {0+sky130_fd_pr__nfet_01v8__eta0_diff_50}
+ etab = -0.043998
+ dsub = 0.45863
* BSIM4 - Sub-threshold parameters
+ voffl = 5.8197729e-9
+ minv = 0.0
* Rout Parameters
+ pclm = {0.12808+sky130_fd_pr__nfet_01v8__pclm_diff_50}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 14.05
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__nfet_01v8__pdits_diff_50}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8__pditsd_diff_50}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.24096074+sky130_fd_pr__nfet_01v8__kt1_diff_50}
+ kt2 = -0.028878939
+ at = 53720.487
+ ute = -1.2690432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.84
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.7
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgso = {2.54e-010*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdl = {0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cf = 1.4067e-12
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.0494e-008+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = {3.6001e-011*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = {2.3347e-010*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.95578
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0.0
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = .2e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8__model.51 nmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 7.39e-07 wmax = 7.41e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__nfet_01v8__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1859e-08+sky130_fd_pr__nfet_01v8__wint_diff}
+ lint = {1.1932e-08+sky130_fd_pr__nfet_01v8__lint_diff}
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.464338660470898+sky130_fd_pr__nfet_01v8__vth0_diff_51+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.127858968273573+sky130_fd_pr__nfet_01v8__k2_diff_51}
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45863
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052000000013
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_51+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__nfet_01v8__nfactor_slope_spectre)
+ nfactor = {2.39756756778143+sky130_fd_pr__nfet_01v8__nfactor_diff_51+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {3.01616370768087e-14+sky130_fd_pr__nfet_01v8__eta0_diff_51}
+ etab = -0.043998
+ u0 = {0.026727469834636+sky130_fd_pr__nfet_01v8__u0_diff_51}
+ ua = {-1.18160361296716e-09+sky130_fd_pr__nfet_01v8__ua_diff_51}
+ ub = {2.07498593195961e-18+sky130_fd_pr__nfet_01v8__ub_diff_51}
+ uc = 7.70039999999991e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {180025.301942316+sky130_fd_pr__nfet_01v8__vsat_diff_51}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_51}
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_51}
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = {0.0+sky130_fd_pr__nfet_01v8__b0_diff_51}
+ b1 = {0.0+sky130_fd_pr__nfet_01v8__b1_diff_51}
+ keta = {-0.0269999999999995+sky130_fd_pr__nfet_01v8__keta_diff_51}
+ dwg = 0.0
+ dwb = 0.0
+ pclm = {0.15158334992144+sky130_fd_pr__nfet_01v8__pclm_diff_51}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__nfet_01v8__pdits_diff_51}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__nfet_01v8__pditsd_diff_51}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_51}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.9999999999999e-8
+ alpha1 = 0.85
+ beta0 = 13.964361997007
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.0494e-08+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ xpart = 0.0
+ cgso = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdo = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ cgdl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgsl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = {3.6001e-11*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = {2.3347e-10*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.236678839850346+sky130_fd_pr__nfet_01v8__kt1_diff_51}
+ kt2 = -0.028878939
+ at = 53720.4869999998
+ ute = -1.29045270074826
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__nfet_01v8__tvoff_diff_51}
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.52 nmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 3.59e-07 wmax = 3.61e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__nfet_01v8__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1859e-08+sky130_fd_pr__nfet_01v8__wint_diff}
+ lint = {1.1932e-08+sky130_fd_pr__nfet_01v8__lint_diff}
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.294216+sky130_fd_pr__nfet_01v8__vth0_diff_52+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.164979+sky130_fd_pr__nfet_01v8__k2_diff_52}
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.745709255106775
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_52+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.11251750684601+sky130_fd_pr__nfet_01v8__nfactor_diff_52}
+ eta0 = {0.0+sky130_fd_pr__nfet_01v8__eta0_diff_52}
+ etab = -0.043998
+ u0 = {0.0420786+sky130_fd_pr__nfet_01v8__u0_diff_52}
+ ua = {-1.21575137545398e-09+sky130_fd_pr__nfet_01v8__ua_diff_52}
+ ub = {3.09344567610299e-18+sky130_fd_pr__nfet_01v8__ub_diff_52}
+ uc = 5.40303933016111e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {205055.7+sky130_fd_pr__nfet_01v8__vsat_diff_52}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_52}
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_52}
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = {0.0+sky130_fd_pr__nfet_01v8__b0_diff_52}
+ b1 = {0.0+sky130_fd_pr__nfet_01v8__b1_diff_52}
+ keta = {-0.140717411247685+sky130_fd_pr__nfet_01v8__keta_diff_52}
+ dwg = 0.0
+ dwb = 0.0
+ pclm = {0.129289552416565+sky130_fd_pr__nfet_01v8__pclm_diff_52}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__nfet_01v8__pdits_diff_52}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__nfet_01v8__pditsd_diff_52}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_52}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.99999998238709e-8
+ alpha1 = 0.85
+ beta0 = 13.8499999988778
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.0494e-08+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ xpart = 0.0
+ cgso = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdo = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ cgdl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgsl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = {3.6001e-11*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = {2.3347e-10*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.240960739938925+sky130_fd_pr__nfet_01v8__kt1_diff_52}
+ kt2 = -0.028878939
+ at = 53720.4870195945
+ ute = -1.19244645977108
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__nfet_01v8__tvoff_diff_52}
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.53 nmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 3.89e-07 wmax = 3.91e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__nfet_01v8__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1859e-08+sky130_fd_pr__nfet_01v8__wint_diff}
+ lint = {1.1932e-08+sky130_fd_pr__nfet_01v8__lint_diff}
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.3288413+sky130_fd_pr__nfet_01v8__vth0_diff_53+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.157868+sky130_fd_pr__nfet_01v8__k2_diff_53}
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.679435816074994
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_53+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.23668316177219+sky130_fd_pr__nfet_01v8__nfactor_diff_53}
+ eta0 = {0.0+sky130_fd_pr__nfet_01v8__eta0_diff_53}
+ etab = -0.043998
+ u0 = {0.0392402+sky130_fd_pr__nfet_01v8__u0_diff_53}
+ ua = {-1.20664055548599e-09+sky130_fd_pr__nfet_01v8__ua_diff_53}
+ ub = {2.8992935911323e-18+sky130_fd_pr__nfet_01v8__ub_diff_53}
+ uc = 6.17577815560697e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {200231.2+sky130_fd_pr__nfet_01v8__vsat_diff_53}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_53}
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_53}
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = {0.0+sky130_fd_pr__nfet_01v8__b0_diff_53}
+ b1 = {0.0+sky130_fd_pr__nfet_01v8__b1_diff_53}
+ keta = {-0.114465726035654+sky130_fd_pr__nfet_01v8__keta_diff_53}
+ dwg = 0.0
+ dwb = 0.0
+ pclm = {0.137157029957607+sky130_fd_pr__nfet_01v8__pclm_diff_53}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__nfet_01v8__pdits_diff_53}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__nfet_01v8__pditsd_diff_53}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_53}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.99999998381496e-8
+ alpha1 = 0.85
+ beta0 = 13.8499999988803
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.0494e-08+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ xpart = 0.0
+ cgso = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdo = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ cgdl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgsl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = {3.6001e-11*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = {2.3347e-10*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.240960739944239+sky130_fd_pr__nfet_01v8__kt1_diff_53}
+ kt2 = -0.028878939
+ at = 53720.4870179085
+ ute = -1.20689692868465
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__nfet_01v8__tvoff_diff_53}
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.54 nmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 5.19e-07 wmax = 5.21e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__nfet_01v8__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1859e-08+sky130_fd_pr__nfet_01v8__wint_diff}
+ lint = {1.1932e-08+sky130_fd_pr__nfet_01v8__lint_diff}
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.418842762400781+sky130_fd_pr__nfet_01v8__vth0_diff_54+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.134449331650343+sky130_fd_pr__nfet_01v8__k2_diff_54}
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.488726498226851
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_54+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.59398387978356+sky130_fd_pr__nfet_01v8__nfactor_diff_54}
+ eta0 = {0.000567585745965331+sky130_fd_pr__nfet_01v8__eta0_diff_54}
+ etab = -0.043998
+ u0 = {0.029403234900804+sky130_fd_pr__nfet_01v8__u0_diff_54}
+ ua = {-1.18042314038701e-09+sky130_fd_pr__nfet_01v8__ua_diff_54}
+ ub = {2.34059900360985e-18+sky130_fd_pr__nfet_01v8__ub_diff_54}
+ uc = 8.3994215401744e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {188589.6289636+sky130_fd_pr__nfet_01v8__vsat_diff_54}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_54}
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_54}
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = {0.0+sky130_fd_pr__nfet_01v8__b0_diff_54}
+ b1 = {0.0+sky130_fd_pr__nfet_01v8__b1_diff_54}
+ keta = {-0.0389235321750072+sky130_fd_pr__nfet_01v8__keta_diff_54}
+ dwg = 0.0
+ dwb = 0.0
+ pclm = {0.15979658657271+sky130_fd_pr__nfet_01v8__pclm_diff_54}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__nfet_01v8__pdits_diff_54}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__nfet_01v8__pditsd_diff_54}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_54}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.99999998792379e-8
+ alpha1 = 0.85
+ beta0 = 13.8499999988876
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.0494e-08+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ xpart = 0.0
+ cgso = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdo = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ cgdl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgsl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = {3.6001e-11*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = {2.3347e-10*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.240960739959532+sky130_fd_pr__nfet_01v8__kt1_diff_54}
+ kt2 = -0.028878939
+ at = 53720.4870130568
+ ute = -1.24847978766035
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__nfet_01v8__tvoff_diff_54}
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.55 nmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 5.39e-07 wmax = 5.41e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__nfet_01v8__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1859e-08+sky130_fd_pr__nfet_01v8__wint_diff}
+ lint = {1.1932e-08+sky130_fd_pr__nfet_01v8__lint_diff}
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.423940356524315+sky130_fd_pr__nfet_01v8__vth0_diff_55+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.133949697045732+sky130_fd_pr__nfet_01v8__k2_diff_55}
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.468254513470327
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_55+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.63233887436463+sky130_fd_pr__nfet_01v8__nfactor_diff_55}
+ eta0 = {0.000653654633574984+sky130_fd_pr__nfet_01v8__eta0_diff_55}
+ etab = -0.043998
+ u0 = {0.029067335067153+sky130_fd_pr__nfet_01v8__u0_diff_55}
+ ua = {-1.17760879167915e-09+sky130_fd_pr__nfet_01v8__ua_diff_55}
+ ub = {2.28062507465678e-18+sky130_fd_pr__nfet_01v8__ub_diff_55}
+ uc = 8.63812195600337e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {187648.696329196+sky130_fd_pr__nfet_01v8__vsat_diff_55}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_55}
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_55}
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = {0.0+sky130_fd_pr__nfet_01v8__b0_diff_55}
+ b1 = {0.0+sky130_fd_pr__nfet_01v8__b1_diff_55}
+ keta = {-0.0308143393015842+sky130_fd_pr__nfet_01v8__keta_diff_55}
+ dwg = 0.0
+ dwb = 0.0
+ pclm = {0.162226864564098+sky130_fd_pr__nfet_01v8__pclm_diff_55}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__nfet_01v8__pdits_diff_55}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__nfet_01v8__pditsd_diff_55}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_55}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.99999998836486e-8
+ alpha1 = 0.85
+ beta0 = 13.8499999988884
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.0494e-08+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ xpart = 0.0
+ cgso = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdo = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ cgdl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgsl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = {3.6001e-11*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = {2.3347e-10*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.240960739961173+sky130_fd_pr__nfet_01v8__kt1_diff_55}
+ kt2 = -0.028878939
+ at = 53720.4870125359
+ ute = -1.25294356355074
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__nfet_01v8__tvoff_diff_55}
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.56 nmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 5.79e-07 wmax = 5.81e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__nfet_01v8__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1859e-08+sky130_fd_pr__nfet_01v8__wint_diff}
+ lint = {1.1932e-08+sky130_fd_pr__nfet_01v8__lint_diff}
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.432023091850352+sky130_fd_pr__nfet_01v8__vth0_diff_56+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.133259025374029+sky130_fd_pr__nfet_01v8__k2_diff_56}
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.458626890941655
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_56+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.58898931986882+sky130_fd_pr__nfet_01v8__nfactor_diff_56}
+ eta0 = {0.000436872496185469+sky130_fd_pr__nfet_01v8__eta0_diff_56}
+ etab = -0.043998
+ u0 = {0.0274613358572528+sky130_fd_pr__nfet_01v8__u0_diff_56}
+ ua = {-1.17807438822708e-09+sky130_fd_pr__nfet_01v8__ua_diff_56}
+ ub = {2.15992684900315e-18+sky130_fd_pr__nfet_01v8__ub_diff_56}
+ uc = 8.36124149707075e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {185147.462677658+sky130_fd_pr__nfet_01v8__vsat_diff_56}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_56}
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_56}
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = {0.0+sky130_fd_pr__nfet_01v8__b0_diff_56}
+ b1 = {0.0+sky130_fd_pr__nfet_01v8__b1_diff_56}
+ keta = {-0.027+sky130_fd_pr__nfet_01v8__keta_diff_56}
+ dwg = 0.0
+ dwb = 0.0
+ pclm = {0.170634292062068+sky130_fd_pr__nfet_01v8__pclm_diff_56}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__nfet_01v8__pdits_diff_56}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__nfet_01v8__pditsd_diff_56}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_56}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.85
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.0494e-08+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ xpart = 0.0
+ cgso = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdo = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ cgdl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgsl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = {3.6001e-11*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = {2.3347e-10*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.2372544684968+sky130_fd_pr__nfet_01v8__kt1_diff_56}
+ kt2 = -0.028878939
+ at = 53720.487
+ ute = -1.27876333778794
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__nfet_01v8__tvoff_diff_56}
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.57 nmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 5.99e-07 wmax = 6.01e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__nfet_01v8__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1859e-08+sky130_fd_pr__nfet_01v8__wint_diff}
+ lint = {1.1932e-08+sky130_fd_pr__nfet_01v8__lint_diff}
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.435490647052556+sky130_fd_pr__nfet_01v8__vth0_diff_57+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.130695574634116+sky130_fd_pr__nfet_01v8__k2_diff_57}
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.458628001829958
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_57+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.55174083029451+sky130_fd_pr__nfet_01v8__nfactor_diff_57}
+ eta0 = {0.000280777222630493+sky130_fd_pr__nfet_01v8__eta0_diff_57}
+ etab = -0.043998
+ u0 = {0.0255723631697938+sky130_fd_pr__nfet_01v8__u0_diff_57}
+ ua = {-1.17916009039874e-09+sky130_fd_pr__nfet_01v8__ua_diff_57}
+ ub = {2.10381012399306e-18+sky130_fd_pr__nfet_01v8__ub_diff_57}
+ uc = 8.12512151367848e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {184781.192020055+sky130_fd_pr__nfet_01v8__vsat_diff_57}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_57}
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_57}
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = {0.0+sky130_fd_pr__nfet_01v8__b0_diff_57}
+ b1 = {0.0+sky130_fd_pr__nfet_01v8__b1_diff_57}
+ keta = {-0.027+sky130_fd_pr__nfet_01v8__keta_diff_57}
+ dwg = 0.0
+ dwb = 0.0
+ pclm = {0.175041865085748+sky130_fd_pr__nfet_01v8__pclm_diff_57}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__nfet_01v8__pdits_diff_57}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__nfet_01v8__pditsd_diff_57}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_57}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.85
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.0494e-08+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ xpart = 0.0
+ cgso = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdo = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ cgdl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgsl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = {3.6001e-11*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = {2.3347e-10*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.235005706750175+sky130_fd_pr__nfet_01v8__kt1_diff_57}
+ kt2 = -0.028878939
+ at = 53720.487
+ ute = -1.29315541296607
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__nfet_01v8__tvoff_diff_57}
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.58 nmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 6.09e-07 wmax = 6.11e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__nfet_01v8__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1859e-08+sky130_fd_pr__nfet_01v8__wint_diff}
+ lint = {1.1932e-08+sky130_fd_pr__nfet_01v8__lint_diff}
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.437287493363183+sky130_fd_pr__nfet_01v8__vth0_diff_58+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.130764442614343+sky130_fd_pr__nfet_01v8__k2_diff_58}
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.458628527848268
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_58+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.53410324470474+sky130_fd_pr__nfet_01v8__nfactor_diff_58}
+ eta0 = {0.000206864326323874+sky130_fd_pr__nfet_01v8__eta0_diff_58}
+ etab = -0.043998
+ u0 = {0.0262837093900552+sky130_fd_pr__nfet_01v8__u0_diff_58}
+ ua = {-1.17967418278736e-09+sky130_fd_pr__nfet_01v8__ua_diff_58}
+ ub = {2.0772382132473e-18+sky130_fd_pr__nfet_01v8__ub_diff_58}
+ uc = 8.01331600252541e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {184824.05082609+sky130_fd_pr__nfet_01v8__vsat_diff_58}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_58}
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_58}
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = {0.0+sky130_fd_pr__nfet_01v8__b0_diff_58}
+ b1 = {0.0+sky130_fd_pr__nfet_01v8__b1_diff_58}
+ keta = {-0.027+sky130_fd_pr__nfet_01v8__keta_diff_58}
+ dwg = 0.0
+ dwb = 0.0
+ pclm = {0.177128901294108+sky130_fd_pr__nfet_01v8__pclm_diff_58}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__nfet_01v8__pdits_diff_58}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__nfet_01v8__pditsd_diff_58}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_58}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.85
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.0494e-08+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ xpart = 0.0
+ cgso = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdo = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ cgdl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgsl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = {3.6001e-11*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = {2.3347e-10*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.233940892358226+sky130_fd_pr__nfet_01v8__kt1_diff_58}
+ kt2 = -0.028878939
+ at = 53720.487
+ ute = -1.29997022507442
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__nfet_01v8__tvoff_diff_58}
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.59 nmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 6.49e-07 wmax = 6.51e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__nfet_01v8__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1859e-08+sky130_fd_pr__nfet_01v8__wint_diff}
+ lint = {1.1932e-08+sky130_fd_pr__nfet_01v8__lint_diff}
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.446590926940662+sky130_fd_pr__nfet_01v8__vth0_diff_59+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.130025900818021+sky130_fd_pr__nfet_01v8__k2_diff_59}
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45863
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.00205199999991097
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_diff_59+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.47472871840281+sky130_fd_pr__nfet_01v8__nfactor_diff_59}
+ eta0 = {3.46392141840565e-15+sky130_fd_pr__nfet_01v8__eta0_diff_59}
+ etab = -0.043998
+ u0 = {0.0283101754480054+sky130_fd_pr__nfet_01v8__u0_diff_59}
+ ua = {-1.18116934445868e-09+sky130_fd_pr__nfet_01v8__ua_diff_59}
+ ub = {2.01115212341674e-18+sky130_fd_pr__nfet_01v8__ub_diff_59}
+ uc = 7.70040000000061e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {179718.751306521+sky130_fd_pr__nfet_01v8__vsat_diff_59}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_59}
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_59}
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = {0.0+sky130_fd_pr__nfet_01v8__b0_diff_59}
+ b1 = {0.0+sky130_fd_pr__nfet_01v8__b1_diff_59}
+ keta = {-0.0270000000000035+sky130_fd_pr__nfet_01v8__keta_diff_59}
+ dwg = 0.0
+ dwb = 0.0
+ pclm = {0.179365413396469+sky130_fd_pr__nfet_01v8__pclm_diff_59}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__nfet_01v8__pdits_diff_59}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__nfet_01v8__pditsd_diff_59}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_59}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0000000000007e-8
+ alpha1 = 0.85
+ beta0 = 13.8631338552423
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.0494e-08+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ xpart = 0.0
+ cgso = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdo = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ cgdl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgsl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = {3.6001e-11*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = {2.3347e-10*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.231617432753867+sky130_fd_pr__nfet_01v8__kt1_diff_59}
+ kt2 = -0.028878939
+ at = 53720.4870000015
+ ute = -1.31575973623066
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__nfet_01v8__tvoff_diff_59}
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.60 nmos
* Model Flag Parameters
+ lmin = 1.79e-07 lmax = 1.81e-07 wmin = 6.49e-07 wmax = 6.51e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__nfet_01v8__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1859e-08+sky130_fd_pr__nfet_01v8__wint_diff}
+ lint = {1.1932e-08+sky130_fd_pr__nfet_01v8__lint_diff}
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.489087926896515+sky130_fd_pr__nfet_01v8__vth0_diff_60+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = {-0.134006560853344+sky130_fd_pr__nfet_01v8__k2_diff_60}
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45863
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.00205200000020338
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.207530000026643+sky130_fd_pr__nfet_01v8__voff_diff_60+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.47472871858988+sky130_fd_pr__nfet_01v8__nfactor_diff_60}
+ eta0 = {2.24339747224379e-10+sky130_fd_pr__nfet_01v8__eta0_diff_60}
+ etab = -0.043998
+ u0 = {0.0290533754484549+sky130_fd_pr__nfet_01v8__u0_diff_60}
+ ua = {-1.18116934443936e-09+sky130_fd_pr__nfet_01v8__ua_diff_60}
+ ub = {2.01115212383615e-18+sky130_fd_pr__nfet_01v8__ub_diff_60}
+ uc = 7.70039999737929e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {186073.551287763+sky130_fd_pr__nfet_01v8__vsat_diff_60}
+ a0 = {1.5+sky130_fd_pr__nfet_01v8__a0_diff_60}
+ ags = {1.25+sky130_fd_pr__nfet_01v8__ags_diff_60}
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = {0.0+sky130_fd_pr__nfet_01v8__b0_diff_60}
+ b1 = {0.0+sky130_fd_pr__nfet_01v8__b1_diff_60}
+ keta = {-0.0270000000140271+sky130_fd_pr__nfet_01v8__keta_diff_60}
+ dwg = 0.0
+ dwb = 0.0
+ pclm = {0.179365413615054+sky130_fd_pr__nfet_01v8__pclm_diff_60}
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__nfet_01v8__pdits_diff_60}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__nfet_01v8__pditsd_diff_60}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_60}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.00000000030811e-8
+ alpha1 = 0.85
+ beta0 = 13.8631338577276
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.0494e-08+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ xpart = 0.0
+ cgso = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdo = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ cgdl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgsl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = {3.6001e-11*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = {2.3347e-10*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.23161743269537+sky130_fd_pr__nfet_01v8__kt1_diff_60}
+ kt2 = -0.028878939
+ at = 53720.4869845596
+ ute = -1.31575973616436
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__nfet_01v8__tvoff_diff_60}
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.61 nmos
* Model Flag Parameters
+ lmin = 2.49e-07 lmax = 2.51e-07 wmin = 6.49e-07 wmax = 6.51e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__nfet_01v8__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1859e-08+sky130_fd_pr__nfet_01v8__wint_diff}
+ lint = {1.1932e-08+sky130_fd_pr__nfet_01v8__lint_diff}
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.516828999955843+sky130_fd_pr__nfet_01v8__vth0_diff_61+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.907073489864784
+ k2 = {-0.141056690055146+sky130_fd_pr__nfet_01v8__k2_diff_61}
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.458630000020494
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.00205199999877256
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.178479999962592+sky130_fd_pr__nfet_01v8__voff_diff_61+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.31430000029416+sky130_fd_pr__nfet_01v8__nfactor_diff_61}
+ eta0 = {0.000694140054006476+sky130_fd_pr__nfet_01v8__eta0_diff_61}
+ etab = -0.0439980000058383
+ u0 = {0.0265683999944639+sky130_fd_pr__nfet_01v8__u0_diff_61}
+ ua = {-1.17321199949531e-09+sky130_fd_pr__nfet_01v8__ua_diff_61}
+ ub = {1.78959100023175e-18+sky130_fd_pr__nfet_01v8__ub_diff_61}
+ uc = 9.25600000175409e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {178031.000033113+sky130_fd_pr__nfet_01v8__vsat_diff_61}
+ a0 = {1.49999999958694+sky130_fd_pr__nfet_01v8__a0_diff_61}
+ ags = {1.24999999991156+sky130_fd_pr__nfet_01v8__ags_diff_61}
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = {0.0+sky130_fd_pr__nfet_01v8__b0_diff_61}
+ b1 = {0.0+sky130_fd_pr__nfet_01v8__b1_diff_61}
+ keta = {-0.08314799998985+sky130_fd_pr__nfet_01v8__keta_diff_61}
+ dwg = 0.0
+ dwb = 0.0
+ pclm = {0.238570000055337+sky130_fd_pr__nfet_01v8__pclm_diff_61}
+ pdiblc1 = 0.356972150070715
+ pdiblc2 = 0.00840611209810397
+ pdiblcb = -0.103295770005614
+ drout = 0.503326659625464
+ pscbe1 = 791419879.962999
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__nfet_01v8__pdits_diff_61}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__nfet_01v8__pditsd_diff_61}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_61}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.16000002175671e-8
+ alpha1 = 0.85
+ beta0 = 14.3199999998433
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.0494e-08+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ xpart = 0.0
+ cgso = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdo = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ cgdl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgsl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = {3.6001e-11*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = {2.3347e-10*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.240960740011289+sky130_fd_pr__nfet_01v8__kt1_diff_61}
+ kt2 = -0.0288789390022443
+ at = 28720.48700069
+ ute = -1.3190431999809
+ ua1 = -2.38473364234619e-11
+ ub1 = 7.07753169398452e-19
+ uc1 = 1.4718625000871e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__nfet_01v8__tvoff_diff_61}
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.62 nmos
* Model Flag Parameters
+ lmin = 4.99e-07 lmax = 5.01e-07 wmin = 6.49e-07 wmax = 6.51e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = {4.148e-09*sky130_fd_pr__nfet_01v8__toxe_mult+MC_MM_SWITCH*GAU*(4.148e-9*sky130_fd_pr__nfet_01v8__toxe_mult*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__nfet_01v8__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1859e-08+sky130_fd_pr__nfet_01v8__wint_diff}
+ lint = {1.1932e-08+sky130_fd_pr__nfet_01v8__lint_diff}
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = {0.565450899957471+sky130_fd_pr__nfet_01v8__vth0_diff_62+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.474984049970259
+ k2 = {-0.011133391990376+sky130_fd_pr__nfet_01v8__k2_diff_62}
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.310307129991228
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = {-0.143636430036188+sky130_fd_pr__nfet_01v8__voff_diff_62+MC_MM_SWITCH*GAU*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.98326009964839+sky130_fd_pr__nfet_01v8__nfactor_diff_62}
+ eta0 = {0.49000000002007+sky130_fd_pr__nfet_01v8__eta0_diff_62}
+ etab = -0.000624999995967518
+ u0 = {0.0229911999984441+sky130_fd_pr__nfet_01v8__u0_diff_62}
+ ua = {-1.4518063001264e-09+sky130_fd_pr__nfet_01v8__ua_diff_62}
+ ub = {1.89644019988929e-18+sky130_fd_pr__nfet_01v8__ub_diff_62}
+ uc = 5.25369999954794e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {186522.999992355+sky130_fd_pr__nfet_01v8__vsat_diff_62}
+ a0 = {1.38460000021864+sky130_fd_pr__nfet_01v8__a0_diff_62}
+ ags = {0.156250000966111+sky130_fd_pr__nfet_01v8__ags_diff_62}
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = {1.82972616194526e-17+sky130_fd_pr__nfet_01v8__b0_diff_62}
+ b1 = {-1.40480910610493e-18+sky130_fd_pr__nfet_01v8__b1_diff_62}
+ keta = {-0.007113313066665+sky130_fd_pr__nfet_01v8__keta_diff_62}
+ dwg = 0.0
+ dwb = 0.0
+ pclm = {0.451809999744611+sky130_fd_pr__nfet_01v8__pclm_diff_62}
+ pdiblc1 = 0.0330317930478704
+ pdiblc2 = 4.64376648463636e-5
+ pdiblcb = -0.0946052099907314
+ drout = 0.999999899967828
+ pscbe1 = 436947010.370449
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__nfet_01v8__pdits_diff_62}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__nfet_01v8__pditsd_diff_62}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {65.968+sky130_fd_pr__nfet_01v8__rdsw_diff_62}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.90000000043483e-6
+ alpha1 = 0.85
+ beta0 = 18.0179999980639
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.0494e-08+sky130_fd_pr__nfet_01v8__dlc_diff+sky130_fd_pr__nfet_01v8__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__nfet_01v8__dwc_diff}
+ xpart = 0.0
+ cgso = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgdo = {2.54e-10*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgbo = 1.0e-13
+ cgdl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ cgsl = {0.0*sky130_fd_pr__nfet_01v8__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = {0.0013459*sky130_fd_pr__nfet_01v8__ajunction_mult}
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = {3.6001e-11*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = {2.3347e-10*sky130_fd_pr__nfet_01v8__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.278949579996893+sky130_fd_pr__nfet_01v8__kt1_diff_62}
+ kt2 = -0.0367185999994936
+ at = 10655.2600384763
+ ute = -1.31027890007953
+ ua1 = 8.3166957016476e-10
+ ub1 = -6.31878999963852e-19
+ uc1 = 5.74042809599642e-12
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__nfet_01v8__tvoff_diff_62}
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
.ends sky130_fd_pr__nfet_01v8
* Well Proximity Effect Parameters
