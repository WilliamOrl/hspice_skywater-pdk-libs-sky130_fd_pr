* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param GAU = AGAUSS(0,1.0,1)
.param sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre = 0.0
* statistics '
*   process '
*   '
*   mismatch '
*     vary sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre dist=gauss std = 1.0
*   '
* '
.subckt  sky130_fd_pr__pfet_g5v0d10v5 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__pfet_g5v0d10v5 d g s b sky130_fd_pr__pfet_g5v0d10v5__model l = 'l' w = 'w' nf = 'nf' ad = 'ad' as = 'as' pd = 'pd' ps = 'ps' nrd = 'nrd' nrs = 'nrs' sa = 'sa' sb = 'sb' sd = 'sd'
.model sky130_fd_pr__pfet_g5v0d10v5__model.0 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.83801+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.9752+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.21432e-8
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.79104
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.1 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.83801+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.9752+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.21432e-8
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.79104
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.2 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.114302440e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.093049466e-7
+ k1 = 6.040731475e-01 lk1 = -6.979374130e-8
+ k2 = 1.794642283e-02 lk2 = 1.928534558e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.968553135e+05 lvsat = -7.626968517e-1
+ ua = 2.452507250e-09 lua = 1.992005672e-15
+ ub = 2.051609960e-19 lub = -2.021653901e-24 wub = -3.673419846e-40 pub = 4.203895393e-45
+ uc = -5.147278145e-11 luc = 9.056405361e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.033771039e-02 lu0 = 4.844372142e-9
+ a0 = 9.137680690e-01 la0 = -1.546789490e-7
+ keta = -4.983044435e-03 lketa = -2.317381043e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.133939896e-01 lags = 1.991943888e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.476254648e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.226775651e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.704496585e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.742918888e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -9.470297320e-03 ltvoff = 7.457480328e-8
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.418324416e-01 lpclm = 5.711948926e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 4.539823206e-03 lpdiblc2 = -1.259176499e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.600987628e+08 lpscbe1 = -1.782698666e+3
+ pscbe2 = -1.504865922e-08 lpscbe2 = 2.366287158e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.790959846e-05 lalpha0 = -2.145230776e-10
+ alpha1 = 0.0
+ beta0 = 3.913253927e+01 lbeta0 = -6.823287865e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.257231195e-08 lagidl = -3.379084961e-15
+ bgidl = 1.480360660e+09 lbgidl = 1.766582567e+3
+ cgidl = 9.305387000e+02 lcgidl = -1.815400047e-3
+ egidl = 1.204746871e+00 legidl = -4.025799642e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.029891654e+00 lkt1 = 1.880861237e-6
+ kt2 = -0.019032
+ at = 6.708935685e+05 lat = -1.896940495e+0
+ ute = -1.222020095e+00 lute = -1.294426000e-6
+ ua1 = 1.369566054e-09 lua1 = -5.220907470e-15
+ ub1 = -2.615148450e-18 lub1 = -4.172369016e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.3 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.407558942e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -9.567978233e-8
+ k1 = 6.022940360e-01 lk1 = -6.290039589e-8
+ k2 = 2.321137301e-02 lk2 = -1.114230396e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.482574000e+04 lvsat = 5.883293380e-2
+ ua = 3.313286986e-09 lua = -1.343171495e-15
+ ub = -1.239166271e-18 lub = 3.574536528e-24
+ uc = -5.443619270e-11 luc = 1.020460868e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.075923934e-02 lu0 = 3.211116053e-9
+ a0 = 8.259928173e-01 la0 = 1.854150415e-7
+ keta = -5.193981200e-03 lketa = -2.235651484e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.379186931e-01 lags = 1.041709726e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-6.458627319e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.046532320e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.228673640e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.469530554e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 1.894059464e-02 ltvoff = -3.550603871e-8
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.020026000e-02 leta0 = 2.317000726e-7
+ etab = -1.214502716e-01 letab = 1.993492223e-7
+ dsub = 8.101185050e-01 ldsub = -9.691091595e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044838468e+00 lpclm = -8.232261816e-7
+ pdiblc1 = 5.780855540e-01 lpdiblc1 = -7.287562876e-7
+ pdiblc2 = -1.089362294e-03 lpdiblc2 = 9.219077146e-9
+ pdiblcb = 1.624600000e-01 lpdiblcb = -7.263325160e-07 wpdiblcb = 2.117582368e-22
+ drout = 1.475880000e-01 ldrout = 1.597931535e-6
+ pscbe1 = -1.515212494e+08 lpscbe1 = 9.745442331e+02 ppscbe1 = 1.734723476e-18
+ pscbe2 = 7.552930057e-08 lpscbe2 = -1.143246472e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.367263259e-05 lalpha0 = -8.186852959e-11
+ alpha1 = -9.373000000e-11 lalpha1 = 3.631662580e-16
+ beta0 = 6.958792439e+01 lbeta0 = -1.248257231e-04 pbeta0 = 4.135903063e-25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.598492210e-09 lagidl = 8.143277003e-15
+ bgidl = 2.607594260e+09 lbgidl = -2.600996740e+3
+ cgidl = 4.558606850e+02 lcgidl = 2.378738990e-5
+ egidl = -1.553543708e+00 legidl = 6.661473036e-06 wegidl = -3.388131789e-21 pegidl = -6.462348536e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -5.065732713e-01 lkt1 = -1.467881698e-7
+ kt2 = -0.019032
+ at = 2.099070230e+05 lat = -1.108020253e-1
+ ute = -1.702412530e+00 lute = 5.669025287e-7
+ ua1 = -4.749579392e-10 lua1 = 1.925885193e-15 wua1 = 7.888609052e-31 pua1 = -2.633107346e-36
+ ub1 = -3.719462890e-18 lub1 = 1.064077136e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.161588576e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 4.567061286e-8
+ k1 = 5.594255100e-01 lk1 = 1.746094295e-8
+ k2 = 1.721982465e-02 lk2 = 1.011752616e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.759635466e+05 lvsat = -1.120139985e-1
+ ua = 3.424749578e-09 lua = -1.552119270e-15
+ ub = 6.432586600e-19 lub = 4.574275196e-26
+ uc = 5.120433160e-13 luc = -9.598764002e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.566702634e-02 lu0 = -5.989021457e-9
+ a0 = 1.000482196e+00 la0 = -1.416827474e-7
+ keta = 4.196097920e-02 lketa = -1.107532036e-07 pketa = 2.019483917e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -2.953636726e-01 lags = 9.164020952e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.577214519e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 6.993797401e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.607583180e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -7.349991292e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.437300000e-05 lcit = -8.197625800e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.695424306e-01 leta0 = -2.357167604e-7
+ etab = -2.832145680e-02 letab = 2.476994612e-8
+ dsub = 7.361665400e-02 ldsub = 4.115372104e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.319675117e-02 lpclm = 9.794673814e-7
+ pdiblc1 = 5.497102520e-03 lpdiblc1 = 3.446180236e-7
+ pdiblc2 = 5.859649450e-03 lpdiblc2 = -3.807540271e-9
+ pdiblcb = -3.999200000e-01 lpdiblcb = 3.279050320e-7
+ drout = 1.515411042e+00 ldrout = -9.661895394e-07 wdrout = 6.776263578e-21
+ pscbe1 = 4.285770285e+08 lpscbe1 = -1.129079987e+2
+ pscbe2 = 1.453315357e-08 lpscbe2 = 1.872993543e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.930920315e-05 lalpha0 = 1.111812197e-10 walpha0 = 6.586988559e-27 palpha0 = -1.825841773e-31
+ alpha1 = 1.874600000e-10 lalpha1 = -1.639525160e-16
+ beta0 = -3.823994821e+01 lbeta0 = 7.730840691e-05 pbeta0 = 5.169878828e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.591291258e-08 lagidl = -3.693735419e-15
+ bgidl = 8.692104800e+08 lbgidl = 6.577774942e+2
+ cgidl = 4.406240220e+02 lcgidl = 5.235003836e-5
+ egidl = 3.067904827e+00 legidl = -2.001894388e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -5.996568654e-01 lkt1 = 2.770633568e-8
+ kt2 = -0.019032
+ at = 2.566266000e+05 lat = -1.983825444e-1
+ ute = -1.219045260e+00 lute = -3.392177556e-7
+ ua1 = 6.683544680e-10 lua1 = -2.173682457e-16
+ ub1 = -3.537019980e-18 lub1 = -2.355997655e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.5 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.569207870e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -6.139003690e-9
+ k1 = 5.897113800e-01 lk1 = -9.027078948e-9
+ k2 = 1.224748260e-02 lk2 = 1.446633652e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.221277900e+04 lvsat = 3.120242289e-2
+ ua = -7.005974442e-10 lua = 2.055909236e-15
+ ub = 3.953608160e-18 lub = -2.849488921e-24 wub = 1.175494351e-38
+ uc = 5.756926820e-12 luc = -5.547051513e-18 puc = 5.877471754e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.034490790e-02 lu0 = -1.334296669e-9
+ a0 = 8.215356750e-01 la0 = 1.482387964e-8
+ keta = -1.503847860e-01 lketa = 5.747240264e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 8.580473760e-01 lags = -9.237120785e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.439968960e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.455676071e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.794710300e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.773260508e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.186500000e-05 lcit = 1.475012900e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -6.676430500e-05 leta0 = 8.344147975e-11
+ etab = 7.176732100e-04 letab = -6.276769895e-10
+ dsub = 1.452643820e+00 ldsub = -7.945599490e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.981899897e+00 lpclm = -6.811383895e-7
+ pdiblc1 = 2.058119406e-01 lpdiblc1 = 1.694226662e-7
+ pdiblc2 = -3.190250770e-02 lpdiblc2 = 2.921924238e-08 ppdiblc2 = -5.048709793e-29
+ pdiblcb = -0.025
+ drout = 3.394990744e-01 ldrout = 6.226306753e-8
+ pscbe1 = -3.957264810e+07 lpscbe1 = 2.965357084e+2
+ pscbe2 = 1.809943684e-08 lpscbe2 = -3.100341415e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.383958563e-04 lalpha0 = -1.491916253e-10
+ alpha1 = 0.0
+ beta0 = 6.636422074e+01 lbeta0 = -1.417839925e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.564856239e-08 lagidl = 4.140193059e-14 pagidl = -9.629649722e-35
+ bgidl = 9.939220000e+08 lbgidl = 5.487047988e+2
+ cgidl = 4.346390400e+02 lcgidl = 5.758450362e-5
+ egidl = 1.783938167e+00 legidl = -8.789371474e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -6.844746740e-01 lkt1 = 1.018879911e-7
+ kt2 = -0.019032
+ at = 4.599040000e+04 lat = -1.416012384e-2
+ ute = -2.035608300e+00 lute = 3.749482792e-7
+ ua1 = -2.737234000e-11 lua1 = 3.911144206e-16
+ ub1 = -4.533281500e-18 lub1 = 6.357305599e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.6 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.616184920e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -7.042993190e-8
+ k1 = 5.931545700e-01 lk1 = -1.134985492e-8
+ k2 = 1.560906540e-02 lk2 = 1.219861276e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.970660440e+04 lvsat = -8.369117282e-4
+ ua = -1.734173913e-09 lua = 2.753159922e-15
+ ub = 2.429225074e-18 lub = -1.821140091e-24 pub = 2.802596929e-45
+ uc = 2.425427600e-12 luc = -3.299622139e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 7.535916100e-03 lu0 = 7.306649199e-9
+ a0 = 9.325686900e-01 la0 = -6.007899227e-8
+ keta = 1.006969500e-02 lketa = -5.077019025e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -5.339122400e-01 lags = 8.466447491e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '5.597797557e-03+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.290154412e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.946105100e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.261914405e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -5.607419160e-02 leta0 = 3.786605193e-08 weta0 = 2.233387654e-23 peta0 = -5.285368065e-29
+ etab = -7.176732100e-04 letab = 3.406077055e-10
+ dsub = 1.951373652e-01 ldsub = 5.375390542e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.727638830e-01 lpclm = 4.718447653e-7
+ pdiblc1 = 1.954452350e-01 lpdiblc1 = 1.764160458e-7
+ pdiblc2 = 2.567465976e-02 lpdiblc2 = -9.622314795e-9
+ pdiblcb = -0.025
+ drout = -6.587081148e-01 ldrout = 7.356536374e-7
+ pscbe1 = 4.300318337e+08 lpscbe1 = -2.025947503e+1
+ pscbe2 = 1.074689378e-08 lpscbe2 = 1.859684134e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.121888374e-04 lalpha0 = 8.731280908e-11 walpha0 = 2.067951531e-25 palpha0 = 9.860761315e-32
+ alpha1 = 0.0
+ beta0 = 2.775061702e+01 lbeta0 = 1.187033782e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.013979700e-08 lagidl = -1.647089666e-14
+ bgidl = 2.044837300e+09 lbgidl = -1.602426626e+2
+ cgidl = 1.208170000e+03 lcgidl = -4.642394820e-4
+ egidl = -1.972262296e-01 legidl = 4.575563545e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -4.343197900e-01 lkt1 = -6.686649367e-8
+ kt2 = -0.019032
+ at = 4.161100000e+04 lat = -1.120578060e-2
+ ute = -1.604382500e+00 lute = 8.404335450e-8
+ ua1 = 5.533492000e-10 lua1 = -6.403303200e-19
+ ub1 = -4.283104100e-18 lub1 = 4.669608859e-25
+ uc1 = -2.698615920e-10 luc1 = 1.083823100e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.7 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.234249940e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -8.855656605e-8
+ k1 = 4.613552000e-01 lk1 = 5.120212608e-8
+ k2 = 3.716517800e-02 lk2 = 1.968081721e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.856701500e+04 lvsat = 9.195937401e-3
+ ua = 1.121182011e-08 lua = -3.391008841e-15
+ ub = -7.305558188e-18 lub = 2.798988045e-24
+ uc = -1.700643000e-12 luc = -1.341389032e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.602169700e-02 lu0 = -6.212702416e-9
+ a0 = 2.303696400e-01 la0 = 2.731846769e-7
+ keta = -1.382421100e-01 lketa = 1.961859241e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.220915536e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 7.699821944e-9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.471062760e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.249936346e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.873000000e-05 lcit = -8.889258000e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.873536240e-01 leta0 = 1.001712706e-7
+ etab = 1.442322380e-02 letab = -6.845262015e-9
+ dsub = 4.160171696e-01 ldsub = -5.107564972e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.006081441e+00 lpclm = 1.238122522e-7
+ pdiblc1 = 1.590305890e+00 lpdiblc1 = -4.855848209e-7
+ pdiblc2 = 7.644681054e-03 lpdiblc2 = -1.065286901e-9
+ pdiblcb = -0.025
+ drout = 8.603890164e-01 ldrout = 1.469013887e-8
+ pscbe1 = 4.798870424e+08 lpscbe1 = -4.392075707e+1
+ pscbe2 = 1.533430865e-08 lpscbe2 = -3.175029615e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.318915270e-05 lalpha0 = 4.507355871e-11
+ alpha1 = 0.0
+ beta0 = 4.555962834e+01 lbeta0 = 3.418181045e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.650368080e-08 lagidl = -5.253195908e-15
+ bgidl = 2.054454200e+09 lbgidl = -1.648068433e+2
+ cgidl = -2.189916000e+03 lcgidl = 1.148492134e-03 wcgidl = -3.469446952e-18 pcgidl = -1.654361225e-24
+ egidl = 1.147431046e+00 legidl = -1.806179887e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -5.000989540e-01 lkt1 = -3.564770243e-8
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.632955400e+00 lute = 9.760405284e-8
+ ua1 = 5.52e-10
+ ub1 = -7.566643200e-18 lub1 = 2.025328543e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.8 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.83801+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.9752+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.21432e-8
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.79104
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.9 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.83801+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.9752+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.21432e-8
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.79104
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.10 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.114302440e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.093049466e-7
+ k1 = 6.040731475e-01 lk1 = -6.979374130e-8
+ k2 = 1.794642283e-02 lk2 = 1.928534558e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.968553135e+05 lvsat = -7.626968517e-1
+ ua = 2.452507250e-09 lua = 1.992005672e-15
+ ub = 2.051609960e-19 lub = -2.021653901e-24 pub = -8.407790786e-45
+ uc = -5.147278145e-11 luc = 9.056405361e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.033771039e-02 lu0 = 4.844372142e-9
+ a0 = 9.137680690e-01 la0 = -1.546789490e-7
+ keta = -4.983044435e-03 lketa = -2.317381043e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.133939896e-01 lags = 1.991943888e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.476254648e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.226775651e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.704496585e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.742918888e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -9.470297320e-03 ltvoff = 7.457480328e-8
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.418324416e-01 lpclm = 5.711948926e-06 wpclm = 1.694065895e-21 ppclm = -6.462348536e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 4.539823206e-03 lpdiblc2 = -1.259176499e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.600987628e+08 lpscbe1 = -1.782698666e+3
+ pscbe2 = -1.504865922e-08 lpscbe2 = 2.366287158e-13 ppscbe2 = 7.703719778e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.790959846e-05 lalpha0 = -2.145230776e-10
+ alpha1 = 0.0
+ beta0 = 3.913253927e+01 lbeta0 = -6.823287865e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.257231195e-08 lagidl = -3.379084961e-15
+ bgidl = 1.480360660e+09 lbgidl = 1.766582567e+3
+ cgidl = 9.305387000e+02 lcgidl = -1.815400047e-3
+ egidl = 1.204746871e+00 legidl = -4.025799642e-06 pegidl = -5.169878828e-26
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.029891654e+00 lkt1 = 1.880861237e-06 wkt1 = 1.355252716e-20
+ kt2 = -0.019032
+ at = 6.708935685e+05 lat = -1.896940495e+0
+ ute = -1.222020095e+00 lute = -1.294426000e-6
+ ua1 = 1.369566054e-09 lua1 = -5.220907470e-15
+ ub1 = -2.615148450e-18 lub1 = -4.172369016e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.11 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.407558942e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -9.567978233e-8
+ k1 = 6.022940360e-01 lk1 = -6.290039589e-8
+ k2 = 2.321137301e-02 lk2 = -1.114230396e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.482574000e+04 lvsat = 5.883293380e-2
+ ua = 3.313286986e-09 lua = -1.343171495e-15
+ ub = -1.239166271e-18 lub = 3.574536528e-24 pub = 1.121038771e-44
+ uc = -5.443619270e-11 luc = 1.020460868e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.075923934e-02 lu0 = 3.211116053e-9
+ a0 = 8.259928173e-01 la0 = 1.854150415e-7
+ keta = -5.193981200e-03 lketa = -2.235651484e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.379186931e-01 lags = 1.041709726e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-6.458627319e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.046532320e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.228673640e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.469530554e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 1.894059464e-02 ltvoff = -3.550603871e-8
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.020026000e-02 leta0 = 2.317000726e-7
+ etab = -1.214502716e-01 letab = 1.993492223e-7
+ dsub = 8.101185050e-01 ldsub = -9.691091595e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044838468e+00 lpclm = -8.232261816e-7
+ pdiblc1 = 5.780855540e-01 lpdiblc1 = -7.287562876e-7
+ pdiblc2 = -1.089362294e-03 lpdiblc2 = 9.219077146e-09 ppdiblc2 = 5.048709793e-29
+ pdiblcb = 1.624600000e-01 lpdiblcb = -7.263325160e-07 wpdiblcb = 8.470329473e-22 ppdiblcb = -1.615587134e-27
+ drout = 1.475880000e-01 ldrout = 1.597931535e-6
+ pscbe1 = -1.515212494e+08 lpscbe1 = 9.745442331e+2
+ pscbe2 = 7.552930057e-08 lpscbe2 = -1.143246472e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.367263259e-05 lalpha0 = -8.186852959e-11
+ alpha1 = -9.373000000e-11 lalpha1 = 3.631662580e-16
+ beta0 = 6.958792439e+01 lbeta0 = -1.248257231e-4
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.598492210e-09 lagidl = 8.143277003e-15
+ bgidl = 2.607594260e+09 lbgidl = -2.600996740e+3
+ cgidl = 4.558606850e+02 lcgidl = 2.378738990e-5
+ egidl = -1.553543708e+00 legidl = 6.661473036e-06 wegidl = 3.388131789e-21
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -5.065732713e-01 lkt1 = -1.467881698e-7
+ kt2 = -0.019032
+ at = 2.099070230e+05 lat = -1.108020253e-1
+ ute = -1.702412530e+00 lute = 5.669025287e-7
+ ua1 = -4.749579392e-10 lua1 = 1.925885193e-15 wua1 = 1.183291358e-30 pua1 = 4.513898307e-36
+ ub1 = -3.719462890e-18 lub1 = 1.064077136e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.12 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.158694739e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 4.512813413e-08 wvth0 = -5.799190771e-09 pvth0 = 1.087116302e-14
+ k1 = 5.594255100e-01 lk1 = 1.746094295e-8
+ k2 = 1.596258392e-02 lk2 = 1.247434964e-08 wk2 = 2.519484790e-08 pk2 = -4.723026188e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.759635466e+05 lvsat = -1.120139985e-01 wvsat = -1.776356839e-15
+ ua = 3.426528736e-09 lua = -1.555454479e-15 wua = -3.565395206e-17 pua = 6.683689852e-23
+ ub = 1.435328217e-18 lub = -1.439070839e-24 wub = -1.587291234e-23 pub = 2.975536147e-29
+ uc = 5.120433160e-13 luc = -9.598764002e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.736949709e-02 lu0 = -9.180473123e-09 wu0 = -3.411716650e-08 pu0 = 6.395604033e-14
+ a0 = 9.873704823e-01 la0 = -1.171035294e-07 wa0 = 2.627560618e-07 pa0 = -4.925625135e-13
+ keta = 4.196097920e-02 lketa = -1.107532036e-7
+ a1 = 0.0
+ a2 = 0.5
+ ags = -3.162150852e-01 lags = 9.554901533e-07 wags = 4.178580550e-07 pags = -7.833167099e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.577214519e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 6.993797401e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.510771171e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.535153370e-07 wnfactor = 1.940092912e-06 pnfactor = -3.636898173e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.437300000e-05 lcit = -8.197625800e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.695778880e-01 leta0 = -2.357832288e-07 weta0 = -7.105590291e-10 peta0 = 1.332013956e-15
+ etab = -2.832145680e-02 letab = 2.476994612e-8
+ dsub = 7.361665400e-02 ldsub = 4.115372104e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.319675117e-02 lpclm = 9.794673814e-7
+ pdiblc1 = 5.497102520e-03 lpdiblc1 = 3.446180236e-7
+ pdiblc2 = 5.859649450e-03 lpdiblc2 = -3.807540271e-9
+ pdiblcb = -3.999200000e-01 lpdiblcb = 3.279050320e-07 ppdiblcb = -3.231174268e-27
+ drout = 1.515411042e+00 ldrout = -9.661895394e-7
+ pscbe1 = 4.285770285e+08 lpscbe1 = -1.129079987e+2
+ pscbe2 = 1.453315357e-08 lpscbe2 = 1.872993543e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.930920315e-05 lalpha0 = 1.111812197e-10 walpha0 = -1.490047809e-25 palpha0 = 1.533596950e-31
+ alpha1 = 1.874600000e-10 lalpha1 = -1.639525160e-16
+ beta0 = -3.823994821e+01 lbeta0 = 7.730840691e-05 wbeta0 = -1.084202172e-19 pbeta0 = -3.618915180e-25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.479575641e-08 lagidl = -2.034551447e-14 wagidl = -1.780103783e-13 pagidl = 3.336982552e-19
+ bgidl = 1.047049931e+09 lbgidl = 3.243996585e+02 wbgidl = -3.563866328e+03 pbgidl = 6.680823819e-3
+ cgidl = 9.210078931e+01 lcgidl = 7.056916904e-04 wcgidl = 6.984334484e-03 pcgidl = -1.309283342e-8
+ egidl = 3.067904827e+00 legidl = -2.001894388e-06 pegidl = -2.584939414e-26
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -5.959711691e-01 lkt1 = 2.079712935e-08 wkt1 = -7.386060245e-08 pkt1 = 1.384590854e-13
+ kt2 = -0.019032
+ at = 2.618881222e+05 lat = -2.082457939e-01 wat = -1.054398322e-01 pat = 1.976575094e-7
+ ute = -1.219045260e+00 lute = -3.392177556e-7
+ ua1 = 6.683544680e-10 lua1 = -2.173682457e-16
+ ub1 = -3.537019980e-18 lub1 = -2.355997655e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.13 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.583677056e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -5.162912393e-09 wvth0 = 2.899595385e-08 pvth0 = -1.956067047e-14
+ k1 = 5.897113800e-01 lk1 = -9.027078948e-9
+ k2 = 1.853368629e-02 lk2 = 1.022566351e-08 wk2 = -1.259742395e-07 pk2 = 8.498222197e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.221277900e+04 lvsat = 3.120242289e-2
+ ua = -7.094932313e-10 lua = 2.061910334e-15 wua = 1.782697603e-16 pua = -1.202607803e-22
+ ub = -6.739624508e-21 lub = -1.778383053e-25 wub = 7.936456169e-23 pub = -5.353933332e-29
+ uc = 5.756926820e-12 luc = -5.547051513e-18 wuc = 2.465190329e-32 puc = -1.175494351e-38
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.183255416e-02 lu0 = 4.408137166e-09 wu0 = 1.705858325e-07 pu0 = -1.150772026e-13
+ a0 = 8.870942420e-01 la0 = -2.940192967e-08 wa0 = -1.313780309e-06 pa0 = 8.862761965e-13
+ keta = -1.503847860e-01 lketa = 5.747240264e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 9.623044390e-01 lags = -1.627030226e-07 wags = -2.089290275e-06 pags = 1.409435219e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.439968960e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.455676071e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '6.278770345e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.099807415e-06 wnfactor = -9.700464562e-06 pnfactor = 6.543933393e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.186500000e-05 lcit = 1.475012900e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -2.440512966e-04 leta0 = 2.030392843e-10 weta0 = 3.552795146e-09 peta0 = -2.396715605e-15
+ etab = 7.176732100e-04 letab = -6.276769895e-10
+ dsub = 1.452643820e+00 ldsub = -7.945599490e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.981899897e+00 lpclm = -6.811383895e-7
+ pdiblc1 = 2.058119406e-01 lpdiblc1 = 1.694226662e-7
+ pdiblc2 = -3.190250770e-02 lpdiblc2 = 2.921924238e-08 wpdiblc2 = 2.117582368e-22 ppdiblc2 = 5.048709793e-29
+ pdiblcb = -0.025
+ drout = 3.394990744e-01 ldrout = 6.226306753e-8
+ pscbe1 = -3.957264810e+07 lpscbe1 = 2.965357084e+2
+ pscbe2 = 1.809943684e-08 lpscbe2 = -3.100341415e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.383958563e-04 lalpha0 = -1.491916253e-10
+ alpha1 = 0.0
+ beta0 = 6.636422074e+01 lbeta0 = -1.417839925e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.006278155e-08 lagidl = 7.136376283e-14 wagidl = 8.900518915e-13 pagidl = -6.004290060e-19
+ bgidl = 1.047247427e+08 lbgidl = 1.148557269e+03 wbgidl = 1.781933164e+04 pbgidl = -1.202092112e-2
+ cgidl = 2.177255203e+03 lcgidl = -1.117984360e-03 wcgidl = -3.492167242e-02 pcgidl = 2.355816022e-8
+ egidl = 1.783938167e+00 legidl = -8.789371474e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -7.029031556e-01 lkt1 = 1.143198448e-07 wkt1 = 3.693030123e-07 pkt1 = -2.491318121e-13
+ kt2 = -0.019032
+ at = 1.968278884e+04 lat = 3.586990651e-03 wat = 5.271991610e-01 pat = -3.556485540e-7
+ ute = -2.035608300e+00 lute = 3.749482792e-7
+ ua1 = -2.737234000e-11 lua1 = 3.911144206e-16
+ ub1 = -4.533281500e-18 lub1 = 6.357305599e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.14 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.616184920e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -7.042993190e-8
+ k1 = 5.931545700e-01 lk1 = -1.134985492e-8
+ k2 = 1.560906540e-02 lk2 = 1.219861276e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.970660440e+04 lvsat = -8.369117282e-4
+ ua = -1.734173913e-09 lua = 2.753159922e-15
+ ub = 2.429225074e-18 lub = -1.821140091e-24 wub = -1.175494351e-38
+ uc = 2.425427600e-12 luc = -3.299622139e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 7.535916100e-03 lu0 = 7.306649199e-9
+ a0 = 9.325686900e-01 la0 = -6.007899227e-8
+ keta = 1.006969500e-02 lketa = -5.077019025e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -5.339122400e-01 lags = 8.466447491e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '5.597797557e-03+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.290154412e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.946105100e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.261914405e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -5.607419160e-02 leta0 = 3.786605193e-08 weta0 = 1.968689858e-22 peta0 = -5.679798518e-29
+ etab = -7.176732100e-04 letab = 3.406077055e-10
+ dsub = 1.951373652e-01 ldsub = 5.375390542e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.727638829e-01 lpclm = 4.718447653e-7
+ pdiblc1 = 1.954452351e-01 lpdiblc1 = 1.764160458e-7
+ pdiblc2 = 2.567465976e-02 lpdiblc2 = -9.622314795e-9
+ pdiblcb = -0.025
+ drout = -6.587081148e-01 ldrout = 7.356536374e-7
+ pscbe1 = 4.300318337e+08 lpscbe1 = -2.025947503e+1
+ pscbe2 = 1.074689378e-08 lpscbe2 = 1.859684134e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.121888374e-04 lalpha0 = 8.731280908e-11 walpha0 = 4.135903063e-25 palpha0 = -3.944304526e-31
+ alpha1 = 0.0
+ beta0 = 2.775061702e+01 lbeta0 = 1.187033782e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.013979700e-08 lagidl = -1.647089666e-14
+ bgidl = 2.044837300e+09 lbgidl = -1.602426626e+2
+ cgidl = 1.208170000e+03 lcgidl = -4.642394820e-4
+ egidl = -1.972262296e-01 legidl = 4.575563545e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -4.343197900e-01 lkt1 = -6.686649367e-8
+ kt2 = -0.019032
+ at = 4.161100000e+04 lat = -1.120578060e-2
+ ute = -1.604382500e+00 lute = 8.404335450e-8
+ ua1 = 5.533492000e-10 lua1 = -6.403303200e-19
+ ub1 = -4.283104100e-18 lub1 = 4.669608859e-25
+ uc1 = -2.698615920e-10 luc1 = 1.083823100e-16 wuc1 = 3.155443621e-30
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.15 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-5.225649209e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.838847567e-07 wvth0 = -4.025194889e-06 pvth0 = 1.910357495e-12
+ k1 = 4.613552000e-01 lk1 = 5.120212608e-8
+ k2 = 6.442202288e-02 lk2 = -1.096801686e-08 wk2 = -5.462216110e-07 pk2 = 2.592367766e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.754295656e+04 lvsat = 4.935955537e-03 wvsat = -1.798760378e-01 pvsat = 8.536916752e-8
+ ua = 1.121022808e-08 lua = -3.390253264e-15 wua = 3.190394850e-17 pua = -1.514161396e-23
+ ub = -5.639724395e-18 lub = 2.008383327e-24 wub = -3.338296940e-23 pub = 1.584355728e-29
+ uc = -1.700643000e-12 luc = -1.341389032e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.018290114e-02 lu0 = -8.187609901e-09 wu0 = -8.338968208e-08 pu0 = 3.957674311e-14
+ a0 = 2.303696400e-01 la0 = 2.731846769e-7
+ keta = -1.382421100e-01 lketa = 1.961859241e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.220915536e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 7.699821944e-9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.209030270e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 2.982242737e-07 wnfactor = 6.537046564e-05 pnfactor = -3.102482299e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.873000000e-05 lcit = -8.889258000e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -3.136432963e-01 leta0 = 1.601083490e-07 weta0 = 2.530819271e-06 peta0 = -1.201126826e-12
+ etab = 1.442322380e-02 letab = -6.845262015e-9
+ dsub = 4.160171696e-01 ldsub = -5.107564972e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.006081441e+00 lpclm = 1.238122522e-7
+ pdiblc1 = 1.590305890e+00 lpdiblc1 = -4.855848209e-7
+ pdiblc2 = 7.644681054e-03 lpdiblc2 = -1.065286901e-9
+ pdiblcb = -0.025
+ drout = 8.603890164e-01 ldrout = 1.469013887e-8
+ pscbe1 = 4.798870424e+08 lpscbe1 = -4.392075707e+1
+ pscbe2 = 1.533430865e-08 lpscbe2 = -3.175029615e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.318915270e-05 lalpha0 = 4.507355871e-11
+ alpha1 = 0.0
+ beta0 = 4.555962834e+01 lbeta0 = 3.418181045e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.693435201e-07 lagidl = -7.304498362e-14 wagidl = -2.862481239e-12 pagidl = 1.358533596e-18
+ bgidl = 2.110793276e+09 lbgidl = -1.915453687e+02 wbgidl = -1.129023586e+03 pbgidl = 5.358345940e-4
+ cgidl = -8.492230377e+03 lcgidl = 4.139570537e-03 wcgidl = 1.262970944e-01 pcgidl = -5.994060102e-8
+ egidl = 1.147431046e+00 legidl = -1.806179887e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -3.319155449e-01 lkt1 = -1.154675484e-07 wkt1 = -3.370361209e-06 pkt1 = 1.599573430e-12
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.632955400e+00 lute = 9.760405284e-8
+ ua1 = 5.52e-10
+ ub1 = -7.566643200e-18 lub1 = 2.025328543e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.16 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.83801+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.9752+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.21432e-8
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.79104
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.17 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.83801+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.9752+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.21432e-8
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.79104
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.18 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.114302440e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.093049466e-7
+ k1 = 6.040731475e-01 lk1 = -6.979374130e-8
+ k2 = 1.794642283e-02 lk2 = 1.928534558e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.968553135e+05 lvsat = -7.626968517e-1
+ ua = 2.452507250e-09 lua = 1.992005672e-15
+ ub = 2.051609960e-19 lub = -2.021653901e-24 pub = 2.802596929e-45
+ uc = -5.147278145e-11 luc = 9.056405361e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.033771038e-02 lu0 = 4.844372142e-9
+ a0 = 9.137680690e-01 la0 = -1.546789490e-7
+ keta = -4.983044435e-03 lketa = -2.317381043e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.133939896e-01 lags = 1.991943888e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.476254648e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.226775651e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.704496585e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.742918888e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -9.470297320e-03 ltvoff = 7.457480328e-8
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.418324416e-01 lpclm = 5.711948926e-06 wpclm = -8.470329473e-22 ppclm = 6.462348536e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 4.539823206e-03 lpdiblc2 = -1.259176499e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.600987628e+08 lpscbe1 = -1.782698666e+3
+ pscbe2 = -1.504865922e-08 lpscbe2 = 2.366287158e-13 ppscbe2 = 3.851859889e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.790959846e-05 lalpha0 = -2.145230776e-10
+ alpha1 = 0.0
+ beta0 = 3.913253927e+01 lbeta0 = -6.823287865e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.257231195e-08 lagidl = -3.379084961e-15
+ bgidl = 1.480360660e+09 lbgidl = 1.766582567e+3
+ cgidl = 9.305387000e+02 lcgidl = -1.815400047e-3
+ egidl = 1.204746871e+00 legidl = -4.025799642e-06 pegidl = -2.584939414e-26
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.029891654e+00 lkt1 = 1.880861237e-6
+ kt2 = -0.019032
+ at = 6.708935685e+05 lat = -1.896940495e+0
+ ute = -1.222020095e+00 lute = -1.294426000e-6
+ ua1 = 1.369566054e-09 lua1 = -5.220907470e-15
+ ub1 = -2.615148450e-18 lub1 = -4.172369016e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.19 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.407558942e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -9.567978233e-8
+ k1 = 6.022940360e-01 lk1 = -6.290039589e-8
+ k2 = 2.321137301e-02 lk2 = -1.114230396e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.482574000e+04 lvsat = 5.883293380e-2
+ ua = 3.313286986e-09 lua = -1.343171495e-15
+ ub = -1.239166271e-18 lub = 3.574536528e-24 pub = -5.605193857e-45
+ uc = -5.443619270e-11 luc = 1.020460868e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.075923934e-02 lu0 = 3.211116053e-9
+ a0 = 8.259928173e-01 la0 = 1.854150415e-7
+ keta = -5.193981200e-03 lketa = -2.235651484e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.379186931e-01 lags = 1.041709726e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-6.458627319e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.046532320e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.228673640e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.469530554e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 1.894059464e-02 ltvoff = -3.550603871e-8
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.020026000e-02 leta0 = 2.317000726e-7
+ etab = -1.214502716e-01 letab = 1.993492223e-7
+ dsub = 8.101185050e-01 ldsub = -9.691091595e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044838468e+00 lpclm = -8.232261816e-7
+ pdiblc1 = 5.780855540e-01 lpdiblc1 = -7.287562876e-7
+ pdiblc2 = -1.089362294e-03 lpdiblc2 = 9.219077146e-09 ppdiblc2 = 2.524354897e-29
+ pdiblcb = 1.624600000e-01 lpdiblcb = -7.263325160e-07 ppdiblcb = -1.615587134e-27
+ drout = 1.475880000e-01 ldrout = 1.597931535e-6
+ pscbe1 = -1.515212494e+08 lpscbe1 = 9.745442331e+02 ppscbe1 = -1.734723476e-18
+ pscbe2 = 7.552930057e-08 lpscbe2 = -1.143246472e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.367263259e-05 lalpha0 = -8.186852959e-11
+ alpha1 = -9.373000000e-11 lalpha1 = 3.631662580e-16
+ beta0 = 6.958792439e+01 lbeta0 = -1.248257231e-4
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.598492210e-09 lagidl = 8.143277003e-15
+ bgidl = 2.607594260e+09 lbgidl = -2.600996740e+3
+ cgidl = 4.558606850e+02 lcgidl = 2.378738990e-5
+ egidl = -1.553543708e+00 legidl = 6.661473036e-06 wegidl = -1.694065895e-21 pegidl = -9.693522803e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -5.065732713e-01 lkt1 = -1.467881698e-7
+ kt2 = -0.019032
+ at = 2.099070230e+05 lat = -1.108020253e-1
+ ute = -1.702412530e+00 lute = 5.669025287e-7
+ ua1 = -4.749579392e-10 lua1 = 1.925885193e-15 wua1 = 5.916456789e-31 pua1 = -2.256949154e-36
+ ub1 = -3.719462890e-18 lub1 = 1.064077136e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.20 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.944259809e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 4.930162240e-09 wvth0 = -3.283049503e-07 pvth0 = 6.154404599e-13
+ k1 = 5.594255100e-01 lk1 = 1.746094295e-8
+ k2 = 1.867375544e-02 lk2 = 7.391987513e-09 wk2 = -1.558061868e-08 pk2 = 2.920742778e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.759635466e+05 lvsat = -1.120139985e-1
+ ua = 3.423722216e-09 lua = -1.550193377e-15 wua = 6.555534084e-18 pua = -1.228900419e-23
+ ub = -2.284352419e-19 lub = 1.679820140e-24 wub = 9.149750675e-24 pub = -1.715212261e-29
+ uc = 5.120433160e-13 luc = -9.598764002e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.186682114e-02 lu0 = 1.134843215e-09 wu0 = 4.864195726e-08 pu0 = -9.118421307e-14
+ a0 = 9.898488547e-01 la0 = -1.217494862e-07 wa0 = 2.254818472e-07 pa0 = -4.226882708e-13
+ keta = 4.196097920e-02 lketa = -1.107532036e-07 pketa = 2.019483917e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -3.137905595e-01 lags = 9.509451374e-07 wags = 3.813936832e-07 pags = -7.149605986e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.577214519e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 6.993797401e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.566712158e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -6.583823106e-07 wnfactor = 1.098751885e-06 pnfactor = -2.059720284e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.437300000e-05 lcit = -8.197625800e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.695306427e-01 leta0 = -2.356946628e-7
+ etab = -2.832145680e-02 letab = 2.476994612e-8
+ dsub = 7.361665400e-02 ldsub = 4.115372104e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.321870319e-02 lpclm = 9.794262302e-07 wpclm = -3.301538117e-10 ppclm = 6.189063353e-16
+ pdiblc1 = 5.497102520e-03 lpdiblc1 = 3.446180236e-7
+ pdiblc2 = 5.859649450e-03 lpdiblc2 = -3.807540271e-9
+ pdiblcb = -3.999200000e-01 lpdiblcb = 3.279050320e-7
+ drout = 1.515411042e+00 ldrout = -9.661895394e-7
+ pscbe1 = 4.285770285e+08 lpscbe1 = -1.129079987e+2
+ pscbe2 = 1.453315357e-08 lpscbe2 = 1.872993543e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.930920315e-05 lalpha0 = 1.111812197e-10 walpha0 = 4.522539570e-26 palpha0 = -1.913614525e-31
+ alpha1 = 1.874600000e-10 lalpha1 = -1.639525160e-16
+ beta0 = -3.823994821e+01 lbeta0 = 7.730840691e-05 wbeta0 = -2.710505431e-20
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.275151873e-08 lagidl = 2.232613486e-15 wagidl = 3.132499365e-15 pagidl = -5.872183310e-21
+ bgidl = 8.100875200e+08 lbgidl = 7.686093950e+2
+ cgidl = 5.564910300e+02 lcgidl = -1.648542548e-4
+ egidl = 3.067904827e+00 legidl = -2.001894388e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -5.771142955e-01 lkt1 = -1.455196595e-08 wkt1 = -3.574641350e-07 pkt1 = 6.701022674e-13
+ kt2 = -0.019032
+ at = 2.517163100e+05 lat = -1.891777147e-01 wat = 4.754214888e-02 pat = -8.912251229e-8
+ ute = -9.624701209e-01 lute = -8.201935114e-07 wute = -3.858837751e-06 pute = 7.233777247e-12
+ ua1 = 9.011863088e-10 lua1 = -6.538348145e-16 wua1 = -3.501743388e-15 pua1 = 6.564368155e-21
+ ub1 = -3.158567259e-18 lub1 = -9.450472355e-25 wub1 = -5.691851713e-24 pub1 = 1.066994522e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.21 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.655851704e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 6.716598934e-08 wvth0 = 1.641524752e-06 pvth0 = -1.107372597e-12
+ k1 = 5.897113800e-01 lk1 = -9.027078948e-9
+ k2 = 4.977828687e-03 lk2 = 1.937044505e-08 wk2 = 7.790309340e-08 pk2 = -5.255342681e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.221277900e+04 lvsat = 3.120242289e-2
+ ua = -6.954606321e-10 lua = 2.052443942e-15 wua = -3.277767042e-17 pua = 2.211181647e-23
+ ub = 8.312077670e-18 lub = -5.789712452e-24 wub = -4.574875337e-23 pub = 3.086210903e-29
+ uc = 5.756926820e-12 luc = -5.547051513e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.934593391e-02 lu0 = -1.415238882e-08 wu0 = -2.432097863e-07 pu0 = 1.640693218e-13
+ a0 = 8.747023803e-01 la0 = -2.104237972e-08 wa0 = -1.127409236e-06 pa0 = 7.605502706e-13
+ keta = -1.503847860e-01 lketa = 5.747240264e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 9.501818106e-01 lags = -1.545250974e-07 wags = -1.906968416e-06 pags = 1.286440894e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.439968960e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.455676071e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.999065412e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.911118467e-06 wnfactor = -5.493759426e-06 pnfactor = 3.706090109e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.186500000e-05 lcit = 1.475012900e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -7.825011000e-06 leta0 = 4.368103202e-11
+ etab = 7.176732100e-04 letab = -6.276769895e-10
+ dsub = 1.452643820e+00 ldsub = -7.945599490e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.981790136e+00 lpclm = -6.810643454e-07 wpclm = 1.650769058e-09 ppclm = -1.113608807e-15
+ pdiblc1 = 2.058119406e-01 lpdiblc1 = 1.694226662e-7
+ pdiblc2 = -3.190250770e-02 lpdiblc2 = 2.921924238e-08 wpdiblc2 = -1.058791184e-22 ppdiblc2 = -2.524354897e-29
+ pdiblcb = -0.025
+ drout = 3.394990744e-01 ldrout = 6.226306753e-8
+ pscbe1 = -3.957264810e+07 lpscbe1 = 2.965357084e+2
+ pscbe2 = 1.809943684e-08 lpscbe2 = -3.100341415e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.383958563e-04 lalpha0 = -1.491916253e-10
+ alpha1 = 0.0
+ beta0 = 6.636422074e+01 lbeta0 = -1.417839925e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.984159316e-08 lagidl = 3.073854914e-14 wagidl = -1.566249683e-14 pagidl = 1.056592036e-20
+ bgidl = 1.289536800e+09 lbgidl = 3.492830547e+2
+ cgidl = -1.446960000e+02 lcgidl = 4.484039216e-4
+ egidl = 1.783938167e+00 legidl = -8.789371474e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -7.971875237e-01 lkt1 = 1.779240795e-07 wkt1 = 1.787320675e-06 pkt1 = -1.205726527e-12
+ kt2 = -0.019032
+ at = 7.054185005e+04 lat = -3.072253204e-02 wat = -2.377107444e-01 pat = 1.603596682e-7
+ ute = -3.318483995e+00 lute = 1.240376223e-06 wute = 1.929418875e-05 pute = -1.301585973e-11
+ ua1 = -1.191531544e-09 lua1 = 1.176456220e-15 wua1 = 1.750871694e-14 pua1 = -1.181138045e-20
+ ub1 = -6.425545103e-18 lub1 = 1.912251586e-24 wub1 = 2.845925856e-23 pub1 = -1.919861583e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.22 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.616184920e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -7.042993190e-8
+ k1 = 5.931545700e-01 lk1 = -1.134985492e-8
+ k2 = 1.560906540e-02 lk2 = 1.219861276e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.970660440e+04 lvsat = -8.369117282e-4
+ ua = -1.734173913e-09 lua = 2.753159922e-15
+ ub = 2.429225074e-18 lub = -1.821140091e-24 wub = 5.877471754e-39 pub = -2.802596929e-45
+ uc = 2.425427600e-12 luc = -3.299622139e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 7.535916100e-03 lu0 = 7.306649199e-9
+ a0 = 9.325686900e-01 la0 = -6.007899227e-8
+ keta = 1.006969500e-02 lketa = -5.077019025e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -5.339122400e-01 lags = 8.466447491e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '5.597797557e-03+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.290154412e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.946105100e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.261914405e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -5.607419160e-02 leta0 = 3.786605193e-08 weta0 = 9.098986738e-24 peta0 = 4.772608477e-29
+ etab = -7.176732100e-04 letab = 3.406077055e-10
+ dsub = 1.951373652e-01 ldsub = 5.375390542e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.727638830e-01 lpclm = 4.718447653e-7
+ pdiblc1 = 1.954452350e-01 lpdiblc1 = 1.764160458e-7
+ pdiblc2 = 2.567465976e-02 lpdiblc2 = -9.622314795e-9
+ pdiblcb = -0.025
+ drout = -6.587081148e-01 ldrout = 7.356536374e-7
+ pscbe1 = 4.300318337e+08 lpscbe1 = -2.025947503e+1
+ pscbe2 = 1.074689378e-08 lpscbe2 = 1.859684134e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.121888374e-04 lalpha0 = 8.731280908e-11 walpha0 = 2.067951531e-25 palpha0 = -9.860761315e-32
+ alpha1 = 0.0
+ beta0 = 2.775061702e+01 lbeta0 = 1.187033782e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.013979700e-08 lagidl = -1.647089666e-14
+ bgidl = 2.044837300e+09 lbgidl = -1.602426626e+2
+ cgidl = 1.208170000e+03 lcgidl = -4.642394820e-04 wcgidl = 6.938893904e-18
+ egidl = -1.972262296e-01 legidl = 4.575563545e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -4.343197900e-01 lkt1 = -6.686649367e-8
+ kt2 = -0.019032
+ at = 4.161100000e+04 lat = -1.120578060e-2
+ ute = -1.604382500e+00 lute = 8.404335450e-8
+ ua1 = 5.533492000e-10 lua1 = -6.403303200e-19
+ ub1 = -4.283104100e-18 lub1 = 4.669608859e-25
+ uc1 = -2.698615920e-10 luc1 = 1.083823100e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.23 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.871047347e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.087416109e-08 wvth0 = 1.457409545e-06 pvth0 = -6.916865699e-13
+ k1 = 4.613552000e-01 lk1 = 5.120212608e-8
+ k2 = 1.658018317e-02 lk2 = 1.173772027e-08 wk2 = 1.733098985e-07 pk2 = -8.225287783e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.906254309e+04 lvsat = 8.960759767e-03 wvsat = -5.233234925e-02 pvsat = 2.483693295e-8
+ ua = 1.120599345e-08 lua = -3.388243508e-15 wua = 9.559194794e-17 pua = -4.536793849e-23
+ ub = -1.014043249e-17 lub = 4.144419391e-24 wub = 3.430676229e-23 pub = -1.628198938e-29
+ uc = -1.700643000e-12 luc = -1.341389032e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.795967952e-02 lu0 = -2.386468919e-09 wu0 = 1.004450776e-07 pu0 = -4.767123383e-14
+ a0 = 2.303696400e-01 la0 = 2.731846769e-7
+ keta = -1.382421100e-01 lketa = 1.961859241e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.220915536e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 7.699821944e-9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '7.613849153e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.266902768e-06 wnfactor = -1.591690778e-05 pnfactor = 7.554164433e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.873000000e-05 lcit = -8.889258000e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.814957342e-01 leta0 = 9.739111607e-08 weta0 = 5.433468946e-07 peta0 = -2.578724362e-13
+ etab = -1.164212229e-02 letab = 5.525351236e-09 wetab = 3.920174878e-07 petab = -1.860514997e-13
+ dsub = 4.160171696e-01 ldsub = -5.107564972e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.019994001e-01 lpclm = 5.054295888e-07 wpclm = 1.209322986e-05 ppclm = -5.739446893e-12
+ pdiblc1 = 1.590305890e+00 lpdiblc1 = -4.855848209e-7
+ pdiblc2 = 7.644681054e-03 lpdiblc2 = -1.065286901e-9
+ pdiblcb = -0.025
+ drout = 8.603890164e-01 ldrout = 1.469013887e-8
+ pscbe1 = 4.798870424e+08 lpscbe1 = -4.392075707e+1
+ pscbe2 = 1.533430865e-08 lpscbe2 = -3.175029615e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.318915270e-05 lalpha0 = 4.507355871e-11
+ alpha1 = 0.0
+ beta0 = 4.555962834e+01 lbeta0 = 3.418181045e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.000559417e-07 lagidl = 5.481200094e-14 wagidl = 1.189231708e-12 pagidl = -5.644093687e-19
+ bgidl = 1.567115115e+09 lbgidl = 6.648428626e+01 wbgidl = 7.047785037e+03 pbgidl = -3.344878779e-3
+ cgidl = -4.873420315e+02 lcgidl = 3.404505282e-04 wcgidl = 5.905206725e-03 pcgidl = -2.802611111e-9
+ egidl = 1.147431046e+00 legidl = -1.806179887e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -7.127423082e-01 lkt1 = 6.527283347e-08 wkt1 = 2.357195622e-06 pkt1 = -1.118725042e-12
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.632955400e+00 lute = 9.760405284e-8
+ ua1 = 5.52e-10
+ ub1 = -7.566643200e-18 lub1 = 2.025328543e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.24 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.83801+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.9752+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.21432e-8
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.79104
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.25 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.83801+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.02039548
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.7054732e-9
+ ub = -5.157e-20
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209529
+ a0 = 0.8941253
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1386898
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.9752+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.21432e-8
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.79104
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.26 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.114302440e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.093049466e-7
+ k1 = 6.040731475e-01 lk1 = -6.979374130e-8
+ k2 = 1.794642283e-02 lk2 = 1.928534558e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.968553135e+05 lvsat = -7.626968517e-1
+ ua = 2.452507250e-09 lua = 1.992005672e-15
+ ub = 2.051609960e-19 lub = -2.021653901e-24 pub = -1.401298464e-45
+ uc = -5.147278145e-11 luc = 9.056405361e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.033771038e-02 lu0 = 4.844372142e-9
+ a0 = 9.137680690e-01 la0 = -1.546789490e-7
+ keta = -4.983044435e-03 lketa = -2.317381043e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.133939896e-01 lags = 1.991943888e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.476254648e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.226775651e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.704496585e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.742918888e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -9.470297320e-03 ltvoff = 7.457480328e-8
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.418324416e-01 lpclm = 5.711948926e-06 wpclm = 8.470329473e-22 ppclm = -6.462348536e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 4.539823206e-03 lpdiblc2 = -1.259176499e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.600987628e+08 lpscbe1 = -1.782698666e+3
+ pscbe2 = -1.504865922e-08 lpscbe2 = 2.366287158e-13 ppscbe2 = -3.851859889e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.790959846e-05 lalpha0 = -2.145230776e-10
+ alpha1 = 0.0
+ beta0 = 3.913253927e+01 lbeta0 = -6.823287865e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.257231195e-08 lagidl = -3.379084961e-15
+ bgidl = 1.480360660e+09 lbgidl = 1.766582567e+3
+ cgidl = 9.305387000e+02 lcgidl = -1.815400047e-3
+ egidl = 1.204746871e+00 legidl = -4.025799642e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.029891654e+00 lkt1 = 1.880861237e-6
+ kt2 = -0.019032
+ at = 6.708935685e+05 lat = -1.896940495e+0
+ ute = -1.222020095e+00 lute = -1.294426000e-6
+ ua1 = 1.369566054e-09 lua1 = -5.220907470e-15
+ ub1 = -2.615148450e-18 lub1 = -4.172369016e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.27 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.407558942e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -9.567978233e-8
+ k1 = 6.022940360e-01 lk1 = -6.290039589e-8
+ k2 = 2.321137301e-02 lk2 = -1.114230396e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.482574000e+04 lvsat = 5.883293380e-2
+ ua = 3.313286986e-09 lua = -1.343171495e-15
+ ub = -1.239166271e-18 lub = 3.574536528e-24 pub = -5.605193857e-45
+ uc = -5.443619270e-11 luc = 1.020460868e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.075923934e-02 lu0 = 3.211116053e-9
+ a0 = 8.259928173e-01 la0 = 1.854150415e-7
+ keta = -5.193981200e-03 lketa = -2.235651484e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.379186931e-01 lags = 1.041709726e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-6.458627319e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.046532320e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.228673640e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.469530554e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 1.894059464e-02 ltvoff = -3.550603871e-8
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.020026000e-02 leta0 = 2.317000726e-7
+ etab = -1.214502716e-01 letab = 1.993492223e-7
+ dsub = 8.101185050e-01 ldsub = -9.691091595e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044838468e+00 lpclm = -8.232261816e-7
+ pdiblc1 = 5.780855540e-01 lpdiblc1 = -7.287562876e-7
+ pdiblc2 = -1.089362294e-03 lpdiblc2 = 9.219077146e-09 ppdiblc2 = 1.262177448e-29
+ pdiblcb = 1.624600000e-01 lpdiblcb = -7.263325160e-07 wpdiblcb = -2.117582368e-22 ppdiblcb = -1.211690350e-27
+ drout = 1.475880000e-01 ldrout = 1.597931535e-6
+ pscbe1 = -1.515212494e+08 lpscbe1 = 9.745442331e+2
+ pscbe2 = 7.552930057e-08 lpscbe2 = -1.143246472e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.367263259e-05 lalpha0 = -8.186852959e-11
+ alpha1 = -9.373000000e-11 lalpha1 = 3.631662580e-16
+ beta0 = 6.958792439e+01 lbeta0 = -1.248257231e-4
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.598492210e-09 lagidl = 8.143277003e-15
+ bgidl = 2.607594260e+09 lbgidl = -2.600996740e+3
+ cgidl = 4.558606850e+02 lcgidl = 2.378738990e-5
+ egidl = -1.553543708e+00 legidl = 6.661473036e-06 wegidl = 8.470329473e-22 pegidl = 1.130910994e-26
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -5.065732713e-01 lkt1 = -1.467881698e-7
+ kt2 = -0.019032
+ at = 2.099070230e+05 lat = -1.108020253e-1
+ ute = -1.702412530e+00 lute = 5.669025287e-7
+ ua1 = -4.749579392e-10 lua1 = 1.925885193e-15 wua1 = -1.972152263e-31 pua1 = -1.880790961e-36
+ ub1 = -3.719462890e-18 lub1 = 1.064077136e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.28 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.271263416e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 6.623025836e-8
+ k1 = 5.594255100e-01 lk1 = 1.746094295e-8
+ k2 = 1.712186945e-02 lk2 = 1.030115298e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.759635466e+05 lvsat = -1.120139985e-1
+ ua = 3.424375171e-09 lua = -1.551417406e-15
+ ub = 6.829130240e-19 lub = -2.859331879e-26
+ uc = 5.120433160e-13 luc = -9.598764002e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.671173604e-02 lu0 = -7.947434261e-9
+ a0 = 1.012307662e+00 la0 = -1.638507671e-7
+ keta = 4.196097920e-02 lketa = -1.107532036e-07 pketa = -1.009741959e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -2.758023690e-01 lags = 8.797324755e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.577214519e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 6.993797401e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.676151820e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -8.635379018e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.437300000e-05 lcit = -8.197625800e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.695306427e-01 leta0 = -2.356946628e-7
+ etab = -2.832145680e-02 letab = 2.476994612e-8
+ dsub = 7.361665400e-02 ldsub = 4.115372104e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.318581867e-02 lpclm = 9.794878755e-7
+ pdiblc1 = 5.497102520e-03 lpdiblc1 = 3.446180236e-7
+ pdiblc2 = 5.859649450e-03 lpdiblc2 = -3.807540271e-9
+ pdiblcb = -3.999200000e-01 lpdiblcb = 3.279050320e-7
+ drout = 1.515411042e+00 ldrout = -9.661895394e-7
+ pscbe1 = 4.285770285e+08 lpscbe1 = -1.129079987e+02 wpscbe1 = 1.818989404e-12
+ pscbe2 = 1.453315357e-08 lpscbe2 = 1.872993543e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.930920315e-05 lalpha0 = 1.111812197e-10 walpha0 = -2.362796183e-26 palpha0 = -8.091538874e-32
+ alpha1 = 1.874600000e-10 lalpha1 = -1.639525160e-16
+ beta0 = -3.823994821e+01 lbeta0 = 7.730840691e-05 pbeta0 = 2.584939414e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.306352700e-08 lagidl = 1.647722786e-15
+ bgidl = 8.100875200e+08 lbgidl = 7.686093950e+2
+ cgidl = 5.564910300e+02 lcgidl = -1.648542548e-4
+ egidl = 3.067904827e+00 legidl = -2.001894388e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -6.127190164e-01 lkt1 = 5.219264394e-8
+ kt2 = -0.019032
+ at = 2.564516800e+05 lat = -1.980546393e-01 wat = 8.881784197e-16
+ ute = -1.346824320e+00 lute = -9.968312973e-8
+ ua1 = 5.524e-10
+ ub1 = -3.725496280e-18 lub1 = 1.177179065e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.29 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.020833670e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -4.313232722e-8
+ k1 = 5.897113800e-01 lk1 = -9.027078948e-9
+ k2 = 1.273725860e-02 lk2 = 1.413593363e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.221277900e+04 lvsat = 3.120242289e-2
+ ua = -6.987254066e-10 lua = 2.054646359e-15
+ ub = 3.755336340e-18 lub = -2.715734751e-24 pub = -5.605193857e-45
+ uc = 5.756926820e-12 luc = -5.547051513e-18 puc = -5.877471754e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.512135940e-02 lu0 = 2.189509149e-9
+ a0 = 7.624083420e-01 la0 = 5.471117849e-8
+ keta = -1.503847860e-01 lketa = 5.747240264e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 7.602408580e-01 lags = -2.639093081e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.439968960e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.455676071e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.451867100e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.541978486e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.186500000e-05 lcit = 1.475012900e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -7.825011000e-06 leta0 = 4.368103202e-11
+ etab = 7.176732100e-04 letab = -6.276769895e-10
+ dsub = 1.452643820e+00 ldsub = -7.945599490e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.981954559e+00 lpclm = -6.811752648e-7
+ pdiblc1 = 2.058119406e-01 lpdiblc1 = 1.694226662e-7
+ pdiblc2 = -3.190250770e-02 lpdiblc2 = 2.921924238e-08 wpdiblc2 = -5.293955920e-23 ppdiblc2 = 1.262177448e-29
+ pdiblcb = -0.025
+ drout = 3.394990744e-01 ldrout = 6.226306753e-8
+ pscbe1 = -3.957264810e+07 lpscbe1 = 2.965357084e+2
+ pscbe2 = 1.809943684e-08 lpscbe2 = -3.100341415e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.383958563e-04 lalpha0 = -1.491916253e-10
+ alpha1 = 0.0
+ beta0 = 6.636422074e+01 lbeta0 = -1.417839925e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.140163450e-08 lagidl = 3.179095303e-14
+ bgidl = 1.289536800e+09 lbgidl = 3.492830547e+2
+ cgidl = -1.446960000e+02 lcgidl = 4.484039216e-4
+ egidl = 1.783938167e+00 legidl = -8.789371474e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -6.191639190e-01 lkt1 = 5.782935576e-8
+ kt2 = -0.019032
+ at = 4.686500000e+04 lat = -1.475012900e-2
+ ute = -1.396713000e+00 lute = -5.605049020e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.30 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.616184920e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -7.042993190e-8
+ k1 = 5.931545700e-01 lk1 = -1.134985492e-8
+ k2 = 1.560906540e-02 lk2 = 1.219861276e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.970660440e+04 lvsat = -8.369117282e-4
+ ua = -1.734173913e-09 lua = 2.753159922e-15
+ ub = 2.429225074e-18 lub = -1.821140091e-24 wub = -2.938735877e-39 pub = 1.401298464e-45
+ uc = 2.425427600e-12 luc = -3.299622139e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 7.535916100e-03 lu0 = 7.306649199e-9
+ a0 = 9.325686900e-01 la0 = -6.007899227e-8
+ keta = 1.006969500e-02 lketa = -5.077019025e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -5.339122400e-01 lags = 8.466447491e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '5.597797557e-03+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.290154412e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.946105100e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.261914405e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -5.607419160e-02 leta0 = 3.786605193e-08 weta0 = -3.226004389e-23 peta0 = 3.194886666e-29
+ etab = -7.176732100e-04 letab = 3.406077055e-10
+ dsub = 1.951373652e-01 ldsub = 5.375390542e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.727638829e-01 lpclm = 4.718447653e-7
+ pdiblc1 = 1.954452350e-01 lpdiblc1 = 1.764160458e-7
+ pdiblc2 = 2.567465976e-02 lpdiblc2 = -9.622314795e-9
+ pdiblcb = -0.025
+ drout = -6.587081148e-01 ldrout = 7.356536374e-7
+ pscbe1 = 4.300318337e+08 lpscbe1 = -2.025947503e+1
+ pscbe2 = 1.074689378e-08 lpscbe2 = 1.859684134e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.121888374e-04 lalpha0 = 8.731280908e-11 walpha0 = 2.067951531e-25 palpha0 = 1.972152263e-31
+ alpha1 = 0.0
+ beta0 = 2.775061702e+01 lbeta0 = 1.187033782e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.013979700e-08 lagidl = -1.647089666e-14
+ bgidl = 2.044837300e+09 lbgidl = -1.602426626e+2
+ cgidl = 1.208170000e+03 lcgidl = -4.642394820e-4
+ egidl = -1.972262296e-01 legidl = 4.575563545e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -4.343197900e-01 lkt1 = -6.686649367e-8
+ kt2 = -0.019032
+ at = 4.161100000e+04 lat = -1.120578060e-2
+ ute = -1.604382500e+00 lute = 8.404335450e-8
+ ua1 = 5.533492000e-10 lua1 = -6.403303200e-19
+ ub1 = -4.283104100e-18 lub1 = 4.669608859e-25
+ uc1 = -2.698615920e-10 luc1 = 1.083823100e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.31 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-5.325902915e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.791267159e-07 wvth0 = -2.101843145e-06 pvth0 = 9.975347566e-13
+ k1 = 4.613552000e-01 lk1 = 5.120212608e-8
+ k2 = 3.578514525e-02 lk2 = 2.623045264e-09 wk2 = -1.950400298e-08 pk2 = 9.256599816e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.903038623e+04 lvsat = 1.846802142e-02 wvsat = 1.487864191e-01 pvsat = -7.061403452e-8
+ ua = 1.122322943e-08 lua = -3.396423707e-15 wua = -7.745383773e-17 pua = 3.675959139e-23
+ ub = -5.634932666e-18 lub = 2.006109172e-24 wub = -1.092753688e-23 pub = 5.186209001e-30
+ uc = -1.700643000e-12 luc = -1.341389032e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.280882728e-02 lu0 = -4.687874446e-09 wu0 = 5.176062330e-08 pu0 = -2.456559182e-14
+ a0 = 2.303696400e-01 la0 = 2.731846769e-7
+ keta = -1.382421100e-01 lketa = 1.961859241e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.220915536e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 7.699821944e-9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '1.102279771e+01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -3.884789751e-06 wnfactor = -5.014205581e-05 pnfactor = 2.379741969e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.873000000e-05 lcit = -8.889258000e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 1.336601363e-02 leta0 = 4.909730531e-09 weta0 = -1.413025302e-06 peta0 = 6.706218084e-13
+ etab = 5.786546728e-02 letab = -2.746295077e-08 wetab = -3.058245318e-07 petab = 1.451443228e-13
+ dsub = 4.160171696e-01 ldsub = -5.107564972e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.346500346e+00 lpclm = -5.123505603e-07 wpclm = -9.437122160e-06 ppclm = 4.478858177e-12
+ pdiblc1 = 1.590305890e+00 lpdiblc1 = -4.855848209e-7
+ pdiblc2 = 7.644681054e-03 lpdiblc2 = -1.065286901e-9
+ pdiblcb = -0.025
+ drout = 8.603890164e-01 ldrout = 1.469013887e-8
+ pscbe1 = 4.798870424e+08 lpscbe1 = -4.392075707e+1
+ pscbe2 = 1.533430865e-08 lpscbe2 = -3.175029615e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.318915270e-05 lalpha0 = 4.507355871e-11
+ alpha1 = 0.0
+ beta0 = 4.555962834e+01 lbeta0 = 3.418181045e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.529197313e-10 lagidl = 6.920655296e-15 wagidl = 1.761273247e-13 pagidl = -8.359002829e-20
+ bgidl = 2.269100000e+09 lbgidl = -2.666777400e+2
+ cgidl = -6.945137266e+02 lcgidl = 4.387742146e-04 wcgidl = 7.985168280e-03 pcgidl = -3.789760866e-9
+ egidl = 1.147431046e+00 legidl = -1.806179887e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -5.629695343e-01 lkt1 = -5.809325017e-09 wkt1 = 8.535075260e-07 pkt1 = -4.050746719e-13
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.632955400e+00 lute = 9.760405284e-8
+ ua1 = 5.52e-10
+ ub1 = -7.566643200e-18 lub1 = 2.025328543e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.32 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.054781168e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = -2.290178211e-7
+ k1 = 0.59521
+ k2 = 2.024960310e-02 wk2 = 1.026943583e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.706056027e-09 wua = -4.102984651e-18
+ ub = 9.722997690e-20 wub = -1.047521482e-24
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.224787558e-02 wu0 = -9.116363924e-9
+ a0 = 8.927673018e-01 wa0 = 9.560030516e-9
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.452740415e-01 wags = -4.635171686e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '6.030281293e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = -7.427557063e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.715843688e-09 wagidl = 3.820748126e-14
+ bgidl = 1704700000.0
+ cgidl = -5.596940000e+01 wcgidl = 5.321870358e-3
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -6.571326203e-01 wkt1 = -9.426806361e-7
+ kt2 = -0.019032
+ at = 3.826259176e+05 wat = 3.335038758e-1
+ ute = -1.009171269e+00 wute = -2.655613309e-6
+ ua1 = 2.431339465e-09 wua1 = -1.214209558e-14
+ ub1 = -1.840448805e-18 wub1 = -9.183774282e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.33 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.054781168e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = -2.290178211e-7
+ k1 = 0.59521
+ k2 = 2.024960310e-02 wk2 = 1.026943583e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.706056027e-09 wua = -4.102984651e-18
+ ub = 9.722997690e-20 wub = -1.047521482e-24
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.224787558e-02 wu0 = -9.116363924e-9
+ a0 = 8.927673018e-01 wa0 = 9.560030516e-9
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.452740415e-01 wags = -4.635171686e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '6.030281293e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = -7.427557063e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.715843688e-09 wagidl = 3.820748126e-14
+ bgidl = 1704700000.0
+ cgidl = -5.596940000e+01 wcgidl = 5.321870358e-3
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -6.571326203e-01 wkt1 = -9.426806361e-7
+ kt2 = -0.019032
+ at = 3.826259176e+05 wat = 3.335038758e-1
+ ute = -1.009171269e+00 wute = -2.655613309e-6
+ ua1 = 2.431339465e-09 wua1 = -1.214209558e-14
+ ub1 = -1.840448805e-18 wub1 = -9.183774282e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.34 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.333023638e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -5.683551847e-07 wvth0 = -5.500043385e-07 pvth0 = 2.527640430e-12
+ k1 = 6.040731475e-01 lk1 = -6.979374130e-8
+ k2 = 1.922459094e-02 lk2 = 8.071560811e-09 wk2 = -8.998042718e-09 pk2 = 7.894275713e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.576337035e+05 lvsat = -1.241302362e+00 wvsat = -4.278674670e-01 pvsat = 3.369285155e-6
+ ua = 2.452255192e-09 lua = 1.998580059e-15 wua = 1.774436570e-18 pua = -4.628234115e-23
+ ub = 2.734357084e-19 lub = -1.387549653e-24 wub = -4.806400470e-25 pub = -4.463964549e-30
+ uc = -5.147278145e-11 luc = 9.056405361e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.141935138e-02 lu0 = 6.524296704e-09 wu0 = -7.614531931e-09 pu0 = -1.182632621e-14
+ a0 = 9.163364768e-01 la0 = -1.855978260e-07 wa0 = -1.808106702e-08 pa0 = 2.176625867e-13
+ keta = -4.983044435e-03 lketa = -2.317381043e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 9.844730333e-02 lags = 3.687418323e-07 wags = 1.052216221e-07 pags = -1.193579415e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.476254648e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.226775651e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '7.768157426e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.368507940e-05 wnfactor = -1.452775133e-05 pnfactor = 5.591118981e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -3.333448060e-02 ltvoff = 2.624957009e-07 wtvoff = 1.679989820e-07 ptvoff = -1.322924783e-12
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.418324416e-01 lpclm = 5.711948926e-06 wpclm = -4.235164736e-22 ppclm = -6.462348536e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 4.539823206e-03 lpdiblc2 = -1.259176499e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.600987628e+08 lpscbe1 = -1.782698666e+3
+ pscbe2 = -1.504865922e-08 lpscbe2 = 2.366287158e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.790959846e-05 lalpha0 = -2.145230776e-10
+ alpha1 = 0.0
+ beta0 = 3.913253927e+01 lbeta0 = -6.823287865e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.832521793e-10 lagidl = 5.826492031e-14 wagidl = 9.331646734e-14 pagidl = -4.339612218e-19
+ bgidl = 1.298513670e+09 lbgidl = 3.198554876e+03 wbgidl = 1.280165714e+03 pbgidl = -1.008079293e-2
+ cgidl = -7.440241817e+01 lcgidl = 1.451526448e-04 wcgidl = 7.074580464e-03 pcgidl = -1.380189100e-8
+ egidl = 1.204746871e+00 legidl = -4.025799642e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.568090750e+00 lkt1 = 7.173430892e-06 wkt1 = 3.788811844e-06 pkt1 = -3.725861069e-11
+ kt2 = -0.019032
+ at = 7.103910885e+05 lat = -2.581019615e+00 wat = -2.780544836e-01 pat = 4.815777457e-6
+ ute = -4.793887545e-01 lute = -4.171825392e-06 wute = -5.227973140e-06 pute = 2.025630473e-11
+ ua1 = 4.765053147e-09 lua1 = -1.837706176e-14 wua1 = -2.390353646e-14 pua1 = 9.261664235e-20
+ ub1 = -4.975337326e-19 lub1 = -1.057491903e-23 wub1 = -1.490757562e-23 pub1 = 4.507264599e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.35 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.872167895e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 2.800164913e-08 wvth0 = 3.270752249e-07 pvth0 = -8.706920465e-13
+ k1 = 6.022940360e-01 lk1 = -6.290039589e-8
+ k2 = 1.899356381e-02 lk2 = 8.966698531e-09 wk2 = 2.969251638e-08 pk2 = -7.096768314e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.311203609e+04 lvsat = 1.951890809e-01 wvsat = 6.894619644e-01 pvsat = -9.599194593e-7
+ ua = 3.316662171e-09 lua = -1.350651224e-15 wua = -2.376061506e-17 pua = 5.265576991e-23
+ ub = -8.095910340e-19 lub = 2.808745763e-24 wub = -3.024122035e-24 pub = 5.391010762e-30
+ uc = -5.443619270e-11 luc = 1.020460868e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.266463995e-02 lu0 = 1.699301589e-09 wu0 = -1.341363161e-08 pu0 = 1.064286541e-14
+ a0 = 8.180318774e-01 la0 = 1.952931749e-07 wa0 = 5.604339259e-08 pa0 = -6.954004453e-14
+ keta = -5.193981200e-03 lketa = -2.235651484e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.765269209e-01 lags = 6.621454604e-08 wags = -2.717940479e-07 pags = 2.672055000e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-6.458627319e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.046532320e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.251479673e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 3.815240221e-06 wnfactor = 6.879246179e-06 pnfactor = -2.703236276e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 6.666896119e-02 ltvoff = -1.249776347e-07 wtvoff = -3.359979639e-07 ptvoff = 6.298617832e-13
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.020026000e-02 leta0 = 2.317000726e-7
+ etab = -1.214502716e-01 letab = 1.993492223e-7
+ dsub = 8.101185050e-01 ldsub = -9.691091595e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044838468e+00 lpclm = -8.232261816e-7
+ pdiblc1 = 5.780855540e-01 lpdiblc1 = -7.287562876e-7
+ pdiblc2 = -1.089362294e-03 lpdiblc2 = 9.219077146e-9
+ pdiblcb = 1.624600000e-01 lpdiblcb = -7.263325160e-07 wpdiblcb = -2.117582368e-22 ppdiblcb = 2.019483917e-28
+ drout = 1.475880000e-01 ldrout = 1.597931535e-6
+ pscbe1 = -1.515212494e+08 lpscbe1 = 9.745442331e+2
+ pscbe2 = 7.552930057e-08 lpscbe2 = -1.143246472e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.367263259e-05 lalpha0 = -8.186852959e-11
+ alpha1 = -9.373000000e-11 lalpha1 = 3.631662580e-16
+ beta0 = 6.958792439e+01 lbeta0 = -1.248257231e-4
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.773065636e-08 lagidl = -1.308160971e-14 wagidl = -5.724877666e-14 pagidl = 1.494188726e-19
+ bgidl = 2.971288240e+09 lbgidl = -3.282777476e+03 wbgidl = -2.560331429e+03 pbgidl = 4.799597297e-3
+ cgidl = -5.107353973e+02 lcgidl = 1.835768406e-03 wcgidl = 6.804639234e-03 pcgidl = -1.275597671e-8
+ egidl = -1.553543708e+00 legidl = 6.661473036e-06 wegidl = 8.470329473e-22 pegidl = 4.846761402e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 5.486180897e-01 lkt1 = -1.027969180e-06 wkt1 = -7.428331922e-06 pkt1 = 6.203334551e-12
+ kt2 = -0.019032
+ at = -1.642614099e+05 lat = 8.079089554e-01 wat = 2.634069437e+00 pat = -6.467537887e-6
+ ute = -1.820035170e+00 lute = 1.022643208e-06 wute = 8.280393884e-07 pute = -3.208321414e-12
+ ua1 = -4.749579392e-10 lua1 = 1.925885193e-15 wua1 = -6.902532921e-31 pua1 = 2.445028250e-36
+ ub1 = -2.648698458e-18 lub1 = -2.240016188e-24 wub1 = -7.537963167e-24 pub1 = 1.651834559e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.36 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.781522521e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.984692673e-07 wvth0 = 3.592120008e-07 pvth0 = -9.309356465e-13
+ k1 = 5.594255100e-01 lk1 = 1.746094295e-8
+ k2 = 9.139407233e-03 lk2 = 2.743930045e-08 wk2 = 5.619490562e-08 pk2 = -1.206490620e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.287255387e+05 lvsat = -7.069963674e-02 wvsat = 3.325459391e-01 pvsat = -2.908446784e-7
+ ua = 3.425946147e-09 lua = -1.555514964e-15 wua = -1.105934828e-17 pua = 2.884597520e-23
+ ub = 2.243229158e-18 lub = -2.914070970e-24 wub = -1.098430728e-23 pub = 2.031317403e-29
+ uc = 5.120433160e-13 luc = -9.598764002e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.199320824e-02 lu0 = -1.578803251e-08 wu0 = -3.718048683e-08 pu0 = 5.519621221e-14
+ a0 = 1.050379372e+00 la0 = -2.402654387e-07 wa0 = -2.680170705e-07 pa0 = 5.379436995e-13
+ keta = 4.196097920e-02 lketa = -1.107532036e-07 pketa = -1.009741959e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.704489964e-01 lags = 7.166556006e-07 wags = -7.416662506e-07 pags = 1.148027931e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-2.251322266e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.963062122e-07 wvoff = 4.745581018e-07 pvoff = -8.896066177e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.845213744e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.046973668e-06 wnfactor = -8.229957454e-06 pnfactor = 1.291350372e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.437300000e-05 lcit = -8.197625800e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.705981493e-01 leta0 = -2.376958107e-07 weta0 = -7.515028683e-09 peta0 = 1.408767277e-14
+ etab = -2.832145680e-02 letab = 2.476994612e-8
+ dsub = -4.667141932e-01 ldsub = 1.424441417e-06 wdsub = 3.803818937e-06 pdsub = -7.130638979e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.318581867e-02 lpclm = 9.794878755e-7
+ pdiblc1 = 5.497102520e-03 lpdiblc1 = 3.446180236e-7
+ pdiblc2 = 5.859649450e-03 lpdiblc2 = -3.807540271e-9
+ pdiblcb = -3.999200000e-01 lpdiblcb = 3.279050320e-07 ppdiblcb = 8.077935669e-28
+ drout = 1.515411042e+00 ldrout = -9.661895394e-7
+ pscbe1 = 4.285770285e+08 lpscbe1 = -1.129079987e+2
+ pscbe2 = 1.453315357e-08 lpscbe2 = 1.872993543e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.930920315e-05 lalpha0 = 1.111812197e-10 walpha0 = -7.113119339e-26 palpha0 = -9.744866976e-32
+ alpha1 = 1.874600000e-10 lalpha1 = -1.639525160e-16
+ beta0 = -3.823994821e+01 lbeta0 = 7.730840691e-05 wbeta0 = -4.065758147e-20
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.133261652e-08 lagidl = 4.140040163e-14 wagidl = 1.717438736e-13 pagidl = -2.798507495e-19
+ bgidl = 5.343792809e+08 lbgidl = 1.285452060e+03 wbgidl = 1.940929759e+03 pbgidl = -3.638466926e-3
+ cgidl = 5.564910300e+02 lcgidl = -1.648542548e-4
+ egidl = 3.067904827e+00 legidl = -2.001894388e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 2.227436344e-02 lkt1 = -4.128523088e-08 wkt1 = -4.470223855e-06 pkt1 = 6.580651692e-13
+ kt2 = -0.019032
+ at = 4.737465164e+05 lat = -3.881007032e-01 wat = -1.529711320e+00 pat = 1.337885520e-6
+ ute = -1.111579041e+00 lute = -3.054286511e-07 wute = -1.656078777e-06 pute = 1.448406498e-12
+ ua1 = 5.524e-10
+ ub1 = -4.064665177e-18 lub1 = 4.143550236e-25 wub1 = 2.387679843e-24 pub1 = -2.088264791e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.37 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-3.301196607e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -3.683000371e-07 wvth0 = -3.322528211e-06 pvth0 = 2.289114343e-12
+ k1 = 5.897113800e-01 lk1 = -9.027078948e-9
+ k2 = 5.825942638e-02 lk2 = -1.552106830e-08 wk2 = -3.204667747e-07 pk2 = 2.087792436e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.829081889e+03 lvsat = 3.416180438e-02 wvsat = 2.382053739e-02 pvsat = -2.083344200e-8
+ ua = -7.199705373e-10 lua = 2.070503768e-15 wua = 1.495613862e-16 pua = -1.116329192e-22
+ ub = -3.921886156e-18 lub = 2.477938884e-24 wub = 5.404608022e-23 pub = -3.656240288e-29
+ uc = 5.756926820e-12 luc = -5.547051513e-18 puc = -5.877471754e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -2.226697881e-03 lu0 = 1.414069738e-08 wu0 = 1.221267843e-07 pu0 = -8.413392708e-14
+ a0 = 5.468225710e-01 la0 = 2.001453396e-07 wa0 = 1.517679848e-06 pa0 = -1.023826826e-12
+ keta = -1.503847860e-01 lketa = 5.747240264e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 4.055667819e-01 lags = 2.128722009e-07 wags = 2.496833142e-06 pags = -1.684363638e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '2.426541837e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -2.128197822e-07 wvoff = -2.372790509e-06 pvoff = 1.600684477e-12
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '8.432400942e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -3.309727592e-06 wnfactor = -2.098235022e-05 pnfactor = 1.244459309e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -2.521241080e-03 ltvoff = 2.205077449e-09 wtvoff = 1.774902287e-08 ptvoff = -1.552329540e-14
+ cit = -1.186500000e-05 lcit = 1.475012900e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.188645822e-04 leta0 = -1.222088285e-09 weta0 = -1.595848491e-09 peta0 = 8.910757774e-15
+ etab = -1.994979222e-03 letab = 1.744808827e-09 wetab = 1.909651974e-08 petab = -1.670181616e-14
+ dsub = 4.154327890e+00 ldsub = -2.617121989e-06 wdsub = -1.901930471e-05 pdsub = 1.283046496e-11
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.981954559e+00 lpclm = -6.811752648e-7
+ pdiblc1 = 2.058119406e-01 lpdiblc1 = 1.694226662e-7
+ pdiblc2 = -3.190250770e-02 lpdiblc2 = 2.921924238e-08 wpdiblc2 = -2.646977960e-23 ppdiblc2 = -3.786532345e-29
+ pdiblcb = -0.025
+ drout = 3.394990744e-01 ldrout = 6.226306753e-8
+ pscbe1 = -3.957264810e+07 lpscbe1 = 2.965357084e+2
+ pscbe2 = 1.809943684e-08 lpscbe2 = -3.100341415e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.383958563e-04 lalpha0 = -1.491916253e-10
+ alpha1 = 0.0
+ beta0 = 6.636422074e+01 lbeta0 = -1.417839925e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.272538524e-08 lagidl = -1.462472671e-14 wagidl = -5.218390971e-13 pagidl = 3.267569166e-19
+ bgidl = 2.668077996e+09 lbgidl = -5.806808359e+02 wbgidl = -9.704648795e+03 pbgidl = 6.546756077e-3
+ cgidl = -1.446960000e+02 lcgidl = 4.484039216e-4
+ egidl = 1.783938167e+00 legidl = -8.789371474e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 9.349458856e-01 lkt1 = -8.395077441e-07 wkt1 = -1.094061599e-05 pkt1 = 6.317070126e-12
+ kt2 = -0.019032
+ at = 4.686500000e+04 lat = -1.475012900e-2
+ ute = -1.396713000e+00 lute = -5.605049020e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.38 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.955234600e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -5.433863406e-08 wvth0 = 2.386840584e-07 pvth0 = -1.132794541e-13
+ k1 = 5.931545700e-01 lk1 = -1.134985492e-8
+ k2 = 2.087032768e-02 lk2 = 9.701617685e-09 wk2 = -3.703821312e-08 pk2 = 1.757833595e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.309030151e+04 lvsat = -2.442814377e-03 wvsat = -2.382053739e-02 pvsat = 1.130522704e-8
+ ua = -1.726546698e-09 lua = 2.749540045e-15 wua = -5.369404027e-17 pua = 2.548319151e-23
+ ub = 2.502321771e-18 lub = -1.855831784e-24 wub = -5.145858366e-25 pub = 2.442224380e-31
+ uc = 2.425427600e-12 luc = -3.299622139e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 8.776860029e-03 lu0 = 6.717697210e-09 wu0 = -8.735992110e-09 pu0 = 4.146101855e-15
+ a0 = 9.325686900e-01 la0 = -6.007899227e-8
+ keta = 1.006969500e-02 lketa = -5.077019025e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -5.339122400e-01 lags = 8.466447491e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '5.597797557e-03+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.290154412e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.160700220e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.102638284e-06 wnfactor = -8.550501866e-06 pnfactor = 4.058068186e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 2.521241080e-03 ltvoff = -1.196581017e-09 wtvoff = -1.774902287e-08 ptvoff = 8.423686256e-15
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -6.163841419e-02 leta0 = 4.050683197e-08 weta0 = 3.917099191e-08 peta0 = -1.859055276e-14
+ etab = 1.994979222e-03 letab = -9.468171386e-10 wetab = -1.909651974e-08 petab = 9.063208268e-15
+ dsub = 1.951075316e-01 ldsub = 5.376806447e-08 wdsub = 2.100228240e-10 pdsub = -9.967683227e-17
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.727638829e-01 lpclm = 4.718447653e-7
+ pdiblc1 = 1.954452350e-01 lpdiblc1 = 1.764160458e-7
+ pdiblc2 = 2.567465976e-02 lpdiblc2 = -9.622314795e-9
+ pdiblcb = -0.025
+ drout = -6.587081148e-01 ldrout = 7.356536374e-7
+ pscbe1 = 4.300318337e+08 lpscbe1 = -2.025947503e+1
+ pscbe2 = 1.074689378e-08 lpscbe2 = 1.859684134e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.121888374e-04 lalpha0 = 8.731280908e-11 walpha0 = -2.067951531e-25 palpha0 = 9.860761315e-32
+ alpha1 = 0.0
+ beta0 = 2.775061702e+01 lbeta0 = 1.187033782e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.809183586e-08 lagidl = -2.499093430e-14 wagidl = -1.263786913e-13 pagidl = 5.997932691e-20
+ bgidl = 2.044837300e+09 lbgidl = -1.602426626e+2
+ cgidl = 1.208170000e+03 lcgidl = -4.642394820e-4
+ egidl = -1.972262296e-01 legidl = 4.575563545e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 3.210070814e-01 lkt1 = -4.253446268e-07 wkt1 = -5.317347088e-06 pkt1 = 2.523612928e-12
+ kt2 = -0.019032
+ at = 4.161100000e+04 lat = -1.120578060e-2
+ ute = -1.604382500e+00 lute = 8.404335450e-8
+ ua1 = 5.533492000e-10 lua1 = -6.403303200e-19
+ ub1 = -4.283104100e-18 lub1 = 4.669608859e-25
+ uc1 = -2.698615920e-10 luc1 = 1.083823100e-16 puc1 = 3.761581923e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.39 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.894478192e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 3.769786678e-08 wvth0 = 1.114340651e-06 pvth0 = -5.288660731e-13
+ k1 = 3.511957926e-01 lk1 = 1.034837808e-07 wk1 = 7.754997555e-07 pk1 = -3.680521840e-13
+ k2 = 1.924232419e-02 lk2 = 1.047426814e-08 wk2 = 9.695408254e-08 pk2 = -4.601440757e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.745021295e+04 lvsat = -1.875002835e-02 wvsat = -4.032731633e-01 pvsat = 1.913934433e-7
+ ua = 1.756642311e-08 lua = -6.406903427e-15 wua = -4.473224333e-14 pua = 2.122992268e-20
+ ub = -6.438912418e-18 lub = 2.387677963e-24 wub = -5.267683429e-24 pub = 2.500042555e-30
+ uc = -4.480346100e-11 luc = 1.911520839e-17 wuc = 3.034350457e-16 puc = -1.440102727e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 6.566136930e-02 lu0 = -2.027969089e-08 wu0 = -1.795145706e-07 pu0 = 8.519761523e-14
+ a0 = -1.287602451e+00 la0 = 9.936142312e-07 wa0 = 1.068621385e-05 pa0 = -5.071677095e-12
+ keta = -4.171339535e-02 lketa = -2.619393557e-08 wketa = -6.795424593e-07 pketa = 3.225108512e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-4.186733391e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.484575373e-07 wvoff = 2.087875267e-06 pvoff = -9.909056018e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.994888515e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -7.474404904e-08 wnfactor = 6.372787194e-06 pnfactor = -3.024524802e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.873000000e-05 lcit = -8.889258000e-12 wcit = 1.033975766e-25
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -5.623675860e-01 leta0 = 2.781528969e-07 weta0 = 2.640021790e-06 peta0 = -1.252954341e-12
+ etab = -4.578875665e-02 letab = 2.173134391e-08 wetab = 4.238800592e-07 petab = -2.011734761e-13
+ dsub = 5.181440022e-01 ldsub = -9.954504447e-08 wdsub = -7.189520677e-07 pdsub = 3.412146513e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.330029082e-01 lpclm = 8.068016844e-07 wpclm = 1.013001373e-05 ppclm = -4.807704518e-12
+ pdiblc1 = 2.521628068e+00 lpdiblc1 = -9.275903269e-07 wpdiblc1 = -6.556318149e-06 ppdiblc1 = 3.111628593e-12
+ pdiblc2 = 3.755248629e-02 lpdiblc2 = -1.525953127e-08 wpdiblc2 = -2.105448477e-07 ppdiblc2 = 9.992458472e-14
+ pdiblcb = -0.025
+ drout = -8.098380068e-01 ldrout = 8.073798841e-07 wdrout = 1.175805752e-05 pdrout = -5.580374098e-12
+ pscbe1 = 5.456931090e+07 lpscbe1 = 1.579350383e+02 wpscbe1 = 2.994150065e+03 ppscbe1 = -1.421023621e-3
+ pscbe2 = 1.507474967e-08 lpscbe2 = -1.943162725e-16 wpscbe2 = 1.827242226e-15 ppscbe2 = -8.672091604e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.239936889e-04 lalpha0 = 2.827553916e-10 walpha0 = 3.525561771e-09 palpha0 = -1.673231616e-15
+ alpha1 = 0.0
+ beta0 = 6.381090558e+00 lbeta0 = 2.201231508e-05 wbeta0 = 2.758089136e-04 pbeta0 = -1.308989104e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.679968219e-07 lagidl = -1.198658407e-13 wagidl = -1.704511249e-12 pagidl = 8.089610389e-19
+ bgidl = 3.350871044e+09 lbgidl = -7.800862776e+02 wbgidl = -7.615447470e+03 pbgidl = 3.614291369e-3
+ cgidl = 2.573111567e+03 lcgidl = -1.112040750e-03 wcgidl = -1.501824719e-02 pcgidl = 7.127660118e-9
+ egidl = 1.232950617e+00 legidl = -2.212055768e-07 wegidl = -6.020403295e-07 pegidl = 2.857283404e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -7.993149162e-02 lkt1 = -2.350591801e-07 wkt1 = -2.546981755e-06 pkt1 = 1.208797541e-12
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.632955400e+00 lute = 9.760405284e-8
+ ua1 = 5.52e-10
+ ub1 = -1.449526402e-17 lub1 = 5.313651986e-24 wub1 = 4.877607717e-23 pub1 = -2.314912622e-29
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.40 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.617872707e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = 5.476882740e-8
+ k1 = 0.59521
+ k2 = 2.024257535e-02 wk2 = 1.062362052e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.705534749e-09 wua = -1.475847549e-18
+ ub = -1.746545158e-20 wub = -4.694799205e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.144958018e-02 wu0 = -5.093117950e-9
+ a0 = 8.923558953e-01 wa0 = 1.163343514e-8
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.501952325e-01 wags = -7.115351577e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.855767916e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = -1.508249247e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -8.997492180e-03 wtvoff = 4.534552510e-8
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.735929641e-09 wagidl = 4.818584415e-14
+ bgidl = 1.596787242e+09 wbgidl = 5.438582861e+2
+ cgidl = 1000.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -9.899838151e-01 wkt1 = 7.348214843e-7
+ kt2 = -0.019032
+ at = 448800.0
+ ute = -1.5361
+ ua1 = 2.2096e-11
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.41 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.617872707e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = 5.476882740e-8
+ k1 = 0.59521
+ k2 = 2.024257535e-02 wk2 = 1.062362052e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.705534749e-09 wua = -1.475847549e-18
+ ub = -1.746545158e-20 wub = -4.694799205e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.144958018e-02 wu0 = -5.093117950e-9
+ a0 = 8.923558953e-01 wa0 = 1.163343514e-8
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.501952325e-01 wags = -7.115351577e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.855767916e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = -1.508249247e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -8.997492180e-03 wtvoff = 4.534552510e-8
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.735929641e-09 wagidl = 4.818584415e-14
+ bgidl = 1.596787242e+09 wbgidl = 5.438582861e+2
+ cgidl = 1000.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -9.899838151e-01 wkt1 = 7.348214843e-7
+ kt2 = -0.019032
+ at = 448800.0
+ ute = -1.5361
+ ua1 = 2.2096e-11
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.42 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.484581968e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.049611250e-07 wvth0 = 3.035756822e-08 pvth0 = 1.922289016e-13
+ k1 = 6.040731475e-01 lk1 = -6.979374130e-8
+ k2 = 1.613894840e-02 lk2 = 3.231442077e-08 wk2 = 6.552966211e-09 pk2 = -4.323631151e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.727359285e+05 lvsat = -5.727663426e-1
+ ua = 2.452535484e-09 lua = 1.992268014e-15 wua = 3.618231383e-19 pua = -1.447092160e-23
+ ub = 3.327024344e-19 lub = -2.757432035e-24 wub = -7.793322559e-25 pub = 2.439963200e-30
+ uc = -5.147278145e-11 luc = 9.056405361e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.112030704e-02 lu0 = 2.592894266e-09 wu0 = -6.107409479e-09 pu0 = 7.987140074e-15
+ a0 = 9.093081526e-01 la0 = -1.334922453e-07 wa0 = 1.734025331e-08 pa0 = -4.493891035e-14
+ keta = -4.983044435e-03 lketa = -2.317381043e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.380856414e-01 lags = 9.535818643e-08 wags = -9.454751549e-08 pags = 1.842183902e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.476254648e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.226775651e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.310106728e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -3.577736407e-06 wnfactor = -2.139677258e-06 pnfactor = 4.972243016e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -1.771291298e-02 ltvoff = 6.863045264e-08 wtvoff = 8.926946799e-08 ptvoff = -3.458834807e-13
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.418324416e-01 lpclm = 5.711948926e-06 wpclm = 2.117582368e-22 ppclm = 3.231174268e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 4.539823206e-03 lpdiblc2 = -1.259176499e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.600987628e+08 lpscbe1 = -1.782698666e+3
+ pscbe2 = -1.504865922e-08 lpscbe2 = 2.366287158e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.790959846e-05 lalpha0 = -2.145230776e-10
+ alpha1 = 0.0
+ beta0 = 3.913253927e+01 lbeta0 = -6.823287865e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.756667635e-10 lagidl = 4.340161705e-14 wagidl = 9.378221799e-14 pagidl = -3.590532054e-19
+ bgidl = 1.340082634e+09 lbgidl = 2.021446106e+03 wbgidl = 1.070666615e+03 pbgidl = -4.148404866e-3
+ cgidl = 1.329341000e+03 lcgidl = -2.593428639e-03 wcgidl = -1.734723476e-18
+ egidl = 1.204746871e+00 legidl = -4.025799642e-06 pegidl = 6.462348536e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.214694827e+00 lkt1 = 1.769509334e-06 wkt1 = 2.007768483e-06 pkt1 = -1.002394843e-11
+ kt2 = -0.019032
+ at = 6.463269298e+05 lat = -1.555445562e+00 wat = 4.481580713e-02 pat = -3.529065548e-7
+ ute = -1.516727000e+00 lute = -1.525546258e-7
+ ua1 = 2.2096e-11
+ ub1 = -3.274419114e-18 lub1 = -3.057556667e-24 wub1 = -9.126397810e-25 pub1 = 7.186673219e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.43 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.930247627e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -3.197435090e-07 wvth0 = -1.476333751e-07 pvth0 = 8.818726105e-13
+ k1 = 6.022940360e-01 lk1 = -6.290039589e-8
+ k2 = 2.850067294e-02 lk2 = -1.558231714e-08 wk2 = -1.822137420e-08 pk2 = 5.275434784e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.379375140e+05 lvsat = -5.047640557e-02 wvsat = -7.179695374e-02 pvsat = 2.781844770e-7
+ ua = 3.313443027e-09 lua = -1.343404356e-15 wua = -7.536786306e-18 pua = 1.613303056e-23
+ ub = -1.427138692e-18 lub = 4.061248394e-24 wub = 8.819218224e-26 pub = -9.213469877e-31
+ uc = -5.443619270e-11 luc = 1.020460868e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.024407360e-02 lu0 = 5.987948356e-09 wu0 = -1.214470988e-09 pu0 = -1.097103940e-14
+ a0 = 8.288190138e-01 la0 = 1.783709719e-07 wa0 = 1.678425714e-09 pa0 = 1.574440684e-14
+ keta = -5.193981200e-03 lketa = -2.235651484e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.272550358e-01 lags = 1.373224510e-07 wags = -2.347379817e-08 pags = -9.116383495e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-6.458627319e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.046532320e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.851847952e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.676766954e-06 wnfactor = -6.226079472e-06 pnfactor = 2.080541703e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.020026000e-02 leta0 = 2.317000726e-7
+ etab = -1.214502716e-01 letab = 1.993492223e-7
+ dsub = 8.101185050e-01 ldsub = -9.691091595e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044837300e+00 lpclm = -8.232216553e-07 wpclm = 5.887350206e-12 ppclm = -2.281112711e-17
+ pdiblc1 = 5.780855540e-01 lpdiblc1 = -7.287562876e-7
+ pdiblc2 = -1.089362294e-03 lpdiblc2 = 9.219077146e-9
+ pdiblcb = 1.624600000e-01 lpdiblcb = -7.263325160e-07 wpdiblcb = -5.293955920e-23
+ drout = 1.475880000e-01 ldrout = 1.597931535e-6
+ pscbe1 = -1.515212494e+08 lpscbe1 = 9.745442331e+2
+ pscbe2 = 7.552930057e-08 lpscbe2 = -1.143246472e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.367263259e-05 lalpha0 = -8.186852959e-11
+ alpha1 = -9.373000000e-11 lalpha1 = 3.631662580e-16
+ beta0 = 6.958792439e+01 lbeta0 = -1.248257231e-4
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.699181308e-08 lagidl = -2.544026035e-14 wagidl = -5.352515725e-14 pagidl = 2.117039507e-19
+ bgidl = 2.463265410e+09 lbgidl = -2.330437878e+03 wbgidl = 3.637978807e-12
+ cgidl = 8.394460850e+02 lcgidl = -6.952818009e-4
+ egidl = -1.553543708e+00 legidl = 6.661473036e-06 wegidl = 4.235164736e-22 pegidl = -1.615587134e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -3.584491878e-01 lkt1 = -1.548100020e-06 wkt1 = -2.856897885e-06 pkt1 = 8.824687876e-12
+ kt2 = -0.019032
+ at = 4.715258448e+05 lat = -8.781612775e-01 wat = -5.701686257e-01 pat = 2.029912128e-6
+ ute = -1.655734990e+00 lute = 3.860457323e-7
+ ua1 = -4.749579392e-10 lua1 = 1.925885193e-15 wua1 = -4.930380658e-32 pua1 = 1.504632769e-36
+ ub1 = -5.262880263e-18 lub1 = 4.646934900e-24 wub1 = 5.636979836e-24 pub1 = -1.819048295e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.665816756e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 5.606279945e-09 wvth0 = 3.008986555e-07 pvth0 = 4.105446597e-14
+ k1 = 5.594255100e-01 lk1 = 1.746094295e-8
+ k2 = 2.297221917e-02 lk2 = -5.218677710e-09 wk2 = -1.351964467e-08 pk2 = 4.394048567e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.662175387e+05 lvsat = -1.034901399e-01 wvsat = 1.435939075e-01 pvsat = -1.255872315e-7
+ ua = 3.420885851e-09 lua = -1.544816673e-15 wua = 1.444350856e-17 pua = -2.507123020e-23
+ ub = -7.542596856e-19 lub = 2.799869408e-24 wub = 4.122425004e-24 pub = -8.483919836e-30
+ uc = 5.120433160e-13 luc = -9.598764002e-19
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.400361766e-02 lu0 = -1.059692941e-09 wu0 = 3.085419786e-09 pu0 = -1.903161465e-14
+ a0 = 9.856332766e-01 la0 = -1.155930452e-07 wa0 = 5.829004264e-08 pa0 = -9.037973025e-14
+ keta = 4.196097920e-02 lketa = -1.107532036e-07 pketa = -2.524354897e-29
+ a1 = 0.0
+ a2 = 0.5
+ ags = -3.856032601e-01 lags = 1.098726612e-06 wags = 3.426673469e-07 pags = -7.775320256e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.031067723e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.643026417e-08 wvoff = -2.049150032e-07 pvoff = 3.841336650e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.392531792e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 8.080671204e-07 wnfactor = 9.170855237e-06 pnfactor = -8.057676772e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 1.509556249e-03 ltvoff = -2.829814145e-09 wtvoff = -7.607855547e-09 ptvoff = 1.426168601e-14
+ cit = 1.437300000e-05 lcit = -8.197625800e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.800716463e-01 leta0 = -2.554548281e-07 weta0 = -5.525952076e-08 peta0 = 1.035894976e-13
+ etab = -2.832145680e-02 letab = 2.476994612e-8
+ dsub = 2.880416713e-01 ldsub = 9.576072890e-09 wdsub = 3.349707444e-12 pdsub = -6.279361574e-18
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.318815502e-02 lpclm = 9.794858321e-07 wpclm = -1.177470041e-11 ppclm = 1.029815298e-17
+ pdiblc1 = 5.497102520e-03 lpdiblc1 = 3.446180236e-7
+ pdiblc2 = 5.859649450e-03 lpdiblc2 = -3.807540271e-9
+ pdiblcb = -3.999200000e-01 lpdiblcb = 3.279050320e-07 wpdiblcb = -4.235164736e-22
+ drout = 1.515411042e+00 ldrout = -9.661895394e-07 wdrout = -1.694065895e-21
+ pscbe1 = 4.285770285e+08 lpscbe1 = -1.129079987e+2
+ pscbe2 = 1.453315357e-08 lpscbe2 = 1.872993543e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.930920315e-05 lalpha0 = 1.111812197e-10 walpha0 = -2.828066345e-28 palpha0 = 1.265922780e-32
+ alpha1 = 1.874600000e-10 lalpha1 = -1.639525160e-16
+ beta0 = -3.823994821e+01 lbeta0 = 7.730840691e-05 wbeta0 = 2.032879073e-20 pbeta0 = -1.938704561e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.076060339e-08 lagidl = -1.375923467e-14 wagidl = 6.039855225e-14 pagidl = -1.857435154e-21
+ bgidl = 9.194999800e+08 lbgidl = 5.635047975e+2
+ cgidl = 1.290266171e+03 lcgidl = -1.540389133e-03 wcgidl = -3.698077018e-03 pcgidl = 6.932415178e-9
+ egidl = 3.067904827e+00 legidl = -2.001894388e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.463015773e+00 lkt1 = 5.225205016e-07 wkt1 = 3.015335435e-06 pkt1 = -2.183400706e-12
+ kt2 = -0.019032
+ at = -2.047692893e+04 lat = 4.414712204e-02 wat = 9.610740228e-01 pat = -8.405553403e-7
+ ute = -1.440179400e+00 lute = -1.803477676e-8
+ ua1 = 5.524e-10
+ ub1 = -2.078259300e-18 lub1 = -1.322955556e-24 wub1 = -7.623400548e-24 pub1 = 6.667426120e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.45 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.291196332e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 2.895142581e-07 wvth0 = 1.521102150e-06 pvth0 = -1.026135511e-12
+ k1 = 5.897113800e-01 lk1 = -9.027078948e-9
+ k2 = -3.719042851e-02 lk2 = 4.739957395e-08 wk2 = 1.605810222e-07 pk2 = -1.083279576e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.355557030e+04 lvsat = 3.002801762e-2
+ ua = -6.779537425e-10 lua = 2.040028436e-15 wua = -6.219468805e-17 pua = 4.195653656e-23
+ ub = 1.164190152e-17 lub = -8.041813179e-24 wub = -2.439223464e-23 pub = 1.645500149e-29
+ uc = 5.756926820e-12 luc = -5.547051513e-18 wuc = -3.081487911e-33 puc = 1.469367939e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.820992232e-02 lu0 = -1.348452700e-08 wu0 = -8.166553251e-08 pu0 = 5.509156823e-14
+ a0 = 8.870498626e-01 la0 = -2.937199129e-08 wa0 = -1.969962948e-07 pa0 = 1.328937005e-13
+ keta = -1.503847860e-01 lketa = 5.747240264e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.375052246e+00 lags = -4.411426929e-07 wags = -2.389175820e-06 pags = 1.611738008e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-4.314535629e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 2.419333036e-07 wvoff = 1.024575016e-06 pvoff = -6.911783057e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.305623527e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -8.651229111e-07 wnfactor = -1.842339094e-07 pnfactor = 1.242841953e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -6.547248256e-03 ltvoff = 4.216667076e-09 wtvoff = 3.803927773e-08 ptvoff = -2.566129676e-14
+ cit = -1.186500000e-05 lcit = 1.475012900e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -5.492095700e-02 leta0 = 3.752970272e-08 weta0 = 2.762976038e-07 peta0 = -1.863903635e-13
+ etab = 1.794166160e-03 letab = -1.569177724e-9
+ dsub = 3.805068940e-01 ldsub = -7.129401086e-08 wdsub = -1.674853722e-11 pdsub = 1.129856321e-17
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.981954559e+00 lpclm = -6.811752648e-7
+ pdiblc1 = 2.058119406e-01 lpdiblc1 = 1.694226662e-7
+ pdiblc2 = -3.190250770e-02 lpdiblc2 = 2.921924238e-08 ppdiblc2 = -6.310887242e-30
+ pdiblcb = -0.025
+ drout = 3.394990744e-01 ldrout = 6.226306753e-8
+ pscbe1 = -3.957264810e+07 lpscbe1 = 2.965357084e+2
+ pscbe2 = 1.809943684e-08 lpscbe2 = -3.100341415e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.383958563e-04 lalpha0 = -1.491916253e-10 palpha0 = 1.972152263e-31
+ alpha1 = 0.0
+ beta0 = 6.636422073e+01 lbeta0 = -1.417839925e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.013829934e-07 lagidl = 8.432155509e-14 wagidl = 2.548356932e-13 pagidl = -1.719121586e-19
+ bgidl = 7.424745000e+08 lbgidl = 7.183312823e+2
+ cgidl = -3.813571703e+03 lcgidl = 2.923427471e-03 wcgidl = 1.849038509e-02 pcgidl = -1.247361378e-8
+ egidl = 1.783938167e+00 legidl = -8.789371474e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.686127331e+00 lkt1 = 7.176538697e-07 wkt1 = 2.269058325e-06 pkt1 = -1.530706746e-12
+ kt2 = -0.019032
+ at = 4.686500000e+04 lat = -1.475012900e-2
+ ute = -1.396713000e+00 lute = -5.605049020e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.46 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-5.566252313e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.060274061e-07 wvth0 = -9.653142790e-07 pvth0 = 6.512010126e-13
+ k1 = 6.187262003e-01 lk1 = -2.860047672e-08 wk1 = -1.288758001e-07 pk1 = 8.693961473e-14
+ k2 = 1.289721619e-02 lk2 = 1.361044884e-08 wk2 = 3.144642230e-09 pk2 = -2.121375648e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.037814089e+05 lvsat = -3.083833313e-02 wvsat = -2.288954178e-01 pvsat = 1.544128489e-7
+ ua = -7.943578928e-09 lua = 6.941419186e-15 wua = 3.127888013e-14 pua = -2.110073253e-20
+ ub = 6.039018427e-18 lub = -4.262108247e-24 wub = -1.833881550e-23 pub = 1.237136493e-29
+ uc = 9.859594647e-12 luc = -8.314711229e-18 wuc = -3.746668535e-17 puc = 2.527502593e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.584765941e-02 lu0 = 2.298271764e-08 wu0 = 1.153665625e-07 pu0 = -7.782628304e-14
+ a0 = 1.067928815e+00 la0 = -1.513929325e-07 wa0 = -6.821874156e-07 pa0 = 4.602036306e-13
+ keta = 2.043996584e-01 lketa = -1.818651835e-07 wketa = -9.793833720e-07 pketa = 6.606920228e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -2.441433232e+00 lags = 2.133458410e-06 wags = 9.613516663e-06 pags = -6.485278341e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '1.247868742e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.333064952e-07 wvoff = -6.006886318e-07 pvoff = 4.052245510e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.388219434e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 4.283578896e-07 wnfactor = 5.422235707e-06 pnfactor = -3.657840208e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -1.000532990e-03 ltvoff = 4.748529571e-10
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.385123935e-01 leta0 = 9.392048579e-08 weta0 = 4.266001655e-07 peta0 = -2.877844716e-13
+ etab = -1.794166160e-03 letab = 8.515112595e-10
+ dsub = 7.403972721e-02 ldsub = 1.354487399e-07 wdsub = 6.103670589e-07 pdsub = -4.117536180e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -7.903108239e-01 lpclm = 1.188994963e-06 wpclm = 5.357679655e-06 ppclm = -3.614290696e-12
+ pdiblc1 = -2.020264446e-01 lpdiblc1 = 4.445504409e-07 wpdiblc1 = 2.003176181e-06 ppdiblc1 = -1.351342652e-12
+ pdiblc2 = 4.735408018e-02 lpdiblc2 = -2.424725181e-08 wpdiblc2 = -1.092598563e-07 ppdiblc2 = 7.370669906e-14
+ pdiblcb = -0.025
+ drout = -2.316162150e+00 ldrout = 1.853772129e-06 wdrout = 8.353230217e-06 pdrout = -5.635089104e-12
+ pscbe1 = 4.756771577e+08 lpscbe1 = -5.105181060e+01 wpscbe1 = -2.300431214e+02 ppscbe1 = 1.551870897e-4
+ pscbe2 = 6.556958714e-09 lpscbe2 = 4.686214331e-15 wpscbe2 = 2.111641799e-14 ppscbe2 = -1.424513558e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.089077284e-04 lalpha0 = 2.200193730e-10 walpha0 = 9.914230801e-10 palpha0 = -6.688140099e-16
+ alpha1 = 0.0
+ beta0 = 1.006320089e+00 lbeta0 = 2.991204053e-05 wbeta0 = 1.347858007e-04 pbeta0 = -9.092650114e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.125640260e-07 lagidl = -6.000710420e-14 wagidl = -3.505094574e-13 pagidl = 2.364536799e-19
+ bgidl = 2.405869767e+09 lbgidl = -4.037951650e+02 wbgidl = -1.819529984e+03 pbgidl = 1.227454927e-3
+ cgidl = 2.254118207e+03 lcgidl = -1.169836142e-03 wcgidl = -5.271365588e-03 pcgidl = 3.556063226e-9
+ egidl = -1.228117110e+00 legidl = 1.152995342e-06 wegidl = 5.195479736e-06 pegidl = -3.504870630e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -4.027877639e-01 lkt1 = -1.480870021e-07 wkt1 = -1.669568722e-06 pkt1 = 1.126291060e-12
+ kt2 = -0.019032
+ at = 4.161100000e+04 lat = -1.120578060e-2
+ ute = -1.712584039e+00 lute = 1.570361125e-07 wute = 5.453136815e-07 pute = -3.678686096e-13
+ ua1 = 5.533492000e-10 lua1 = -6.403303200e-19
+ ub1 = -4.283104100e-18 lub1 = 4.669608859e-25
+ uc1 = -2.698615920e-10 luc1 = 1.083823100e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.47 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.014532223e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.129525208e-08 wvth0 = 1.240760929e-06 pvth0 = -3.958022811e-13
+ k1 = 3.535506861e-01 lk1 = 9.725182232e-08 wk1 = 7.636315727e-07 pk1 = -3.366443844e-13
+ k2 = 8.119398500e-02 lk2 = -1.880319764e-08 wk2 = -2.152696498e-07 pk2 = 1.015380473e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.431817254e+05 lvsat = -4.953772330e-02 wvsat = -6.337506567e-01 pvsat = 3.465571452e-7
+ ua = 1.976349271e-08 lua = -6.208357013e-15 wua = -5.580502589e-14 pua = 2.022928926e-20
+ ub = -1.627171550e-17 lub = 6.326566076e-24 wub = 4.428763822e-23 pub = -1.735115000e-29
+ uc = -1.483631033e-10 luc = 6.677778123e-17 wuc = 8.253545169e-16 puc = -3.842199166e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 6.086328266e-02 lu0 = -1.342429547e-08 wu0 = -1.553331928e-07 pu0 = 5.064782079e-14
+ a0 = 1.284724417e+00 la0 = -2.542841253e-07 wa0 = -2.277788806e-06 pa0 = 1.217476050e-12
+ keta = -1.396567566e-01 lketa = -1.857600899e-08 wketa = -1.859278990e-07 pketa = 2.841180553e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -9.701081995e-01 lags = 1.435167550e-06 wags = 1.118889242e-05 pags = -7.232951677e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.713618190e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 7.245674543e-09 wvoff = 8.414756572e-07 pvoff = -2.792266205e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.138643809e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -8.769935186e-07 wnfactor = -4.431302163e-06 pnfactor = 1.018648865e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.719768954e-05 lcit = -2.240002346e-11 wcit = -1.434713479e-10 pcit = 6.809150170e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 7.198875442e-01 leta0 = -3.134761247e-07 weta0 = -3.822282487e-06 peta0 = 1.728735235e-12
+ etab = 1.053906255e-02 letab = -5.001839085e-09 wetab = 1.399993413e-07 petab = -6.644368736e-14
+ dsub = 6.328581824e-01 ldsub = -1.297664990e-07 wdsub = -1.297088135e-06 pdsub = 4.935246168e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.094281559e-01 lpclm = 6.195988427e-07 wpclm = 5.884333027e-06 ppclm = -3.864240386e-12
+ pdiblc1 = 8.578265186e-01 lpdiblc1 = -5.845577546e-08 wpdiblc1 = 1.828902246e-06 ppdiblc1 = -1.268632242e-12
+ pdiblc2 = -7.115810279e-02 lpdiblc2 = 3.199863023e-08 wpdiblc2 = 3.373343443e-07 ppdiblc2 = -1.382469086e-13
+ pdiblcb = -1.163707582e+00 lpdiblcb = 5.404306182e-07 wpdiblcb = 5.738853915e-06 ppdiblcb = -2.723660068e-12
+ drout = 6.417129410e+00 ldrout = -2.291048045e-06 wdrout = -2.466438396e-05 pdrout = 1.003507059e-11
+ pscbe1 = 8.464049832e+08 lpscbe1 = -2.269992366e+02 wpscbe1 = -9.965401889e+02 ppscbe1 = 5.189665979e-4
+ pscbe2 = 2.429493870e-08 lpscbe2 = -3.732230970e-15 wpscbe2 = -4.464062953e-14 ppscbe2 = 1.696315918e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.180099375e-04 lalpha0 = -7.751575129e-11 walpha0 = -7.179647375e-10 palpha0 = 1.424614484e-16
+ alpha1 = 5.693537908e-10 lalpha1 = -2.702153091e-16 walpha1 = -2.869426957e-15 palpha1 = 1.361830034e-21
+ beta0 = -1.560409627e+02 lbeta0 = 1.044466809e-04 wbeta0 = 1.094382928e-03 pbeta0 = -5.463512976e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.382644799e-07 lagidl = -1.196645396e-13 wagidl = -1.554666311e-12 pagidl = 8.079465226e-19
+ bgidl = -1.454027607e+09 lbgidl = 1.428112129e+03 wbgidl = 1.660026153e+04 pbgidl = -7.514578128e-3
+ cgidl = -4.011031773e+02 lcgidl = 9.033192659e-05 wcgidl = -2.881162040e-05 pcgidl = 1.067947113e-9
+ egidl = 1.072303609e+01 legidl = -4.519021967e-06 wegidl = -4.843013515e-05 pegidl = 2.194584619e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.223343184e+00 lkt1 = 2.413486003e-07 wkt1 = 3.215579918e-06 pkt1 = -1.192200485e-12
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -8.471985320e-01 lute = -2.536758490e-07 wute = -3.960054321e-06 pute = 1.770379044e-12
+ ua1 = 5.52e-10
+ ub1 = -4.817079200e-18 lub1 = 7.203854683e-25
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.48 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.799141448e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = 1.098708267e-7
+ k1 = 6.093966538e-01 wk1 = -4.312453352e-8
+ k2 = 1.296940685e-01 wk2 = -3.316478489e-7
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.201713276e+05 wvsat = -6.131672095e-2
+ ua = 2.730945098e-09 wua = -7.871812552e-17
+ ub = -1.494700396e-19 wub = -6.821290178e-26
+ uc = -5.673011313e-11 wuc = 5.094124527e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.033951309e-02 wu0 = -1.718740453e-9
+ a0 = 8.300474084e-01 wa0 = 2.010385245e-7
+ keta = -6.186135826e-03 wketa = -5.288528177e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.182081156e-01 wags = 2.608079422e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-8.724108458e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' wvoff = -1.812804359e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.054823045e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = 9.264597685e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 9.050615880e-03 wtvoff = -9.517041590e-9
+ cit = 1.513265333e-05 wcit = -1.560221907e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.947442565e-01 wpclm = 2.365798772e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 4.635371898e-03 wpdiblc2 = -5.151190267e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 4.521724980e+08 wpscbe1 = -3.600932249e+2
+ pscbe2 = 1.501717205e-08 wpscbe2 = -4.928741005e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.199314476e-05 walpha0 = -9.522451503e-11
+ alpha1 = 0.0
+ beta0 = 3.908397742e+01 wbeta0 = -2.486344668e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.807909118e-09 wagidl = 3.884765322e-14
+ bgidl = 1.758248979e+09 wbgidl = 5.304754484e+1
+ cgidl = 1.546114315e+03 wcgidl = -1.660076109e-3
+ egidl = 4.898457770e-01 wegidl = 6.190923707e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -7.715522461e-01 wkt1 = 7.083407459e-8
+ kt2 = -0.019032
+ at = 5.588748834e+05 wat = -3.346051902e-1
+ ute = -1.515569387e+00 wute = -6.240887629e-8
+ ua1 = 2.2096e-11
+ ub1 = -3.569388362e-18 wub1 = -2.836483427e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.49 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.799141448e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = 1.098708267e-7
+ k1 = 6.093966538e-01 wk1 = -4.312453352e-8
+ k2 = 1.296940685e-01 wk2 = -3.316478489e-7
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.201713276e+05 wvsat = -6.131672095e-2
+ ua = 2.730945098e-09 wua = -7.871812552e-17
+ ub = -1.494700396e-19 wub = -6.821290178e-26
+ uc = -5.673011313e-11 wuc = 5.094124527e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.033951309e-02 wu0 = -1.718740453e-9
+ a0 = 8.300474084e-01 wa0 = 2.010385245e-7
+ keta = -6.186135826e-03 wketa = -5.288528177e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.182081156e-01 wags = 2.608079422e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-8.724108458e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' wvoff = -1.812804359e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.054823045e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = 9.264597685e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 9.050615880e-03 wtvoff = -9.517041590e-9
+ cit = 1.513265333e-05 wcit = -1.560221907e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.947442565e-01 wpclm = 2.365798772e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 4.635371898e-03 wpdiblc2 = -5.151190267e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 4.521724980e+08 wpscbe1 = -3.600932249e+2
+ pscbe2 = 1.501717205e-08 wpscbe2 = -4.928741005e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.199314476e-05 walpha0 = -9.522451503e-11
+ alpha1 = 0.0
+ beta0 = 3.908397742e+01 wbeta0 = -2.486344668e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.807909118e-09 wagidl = 3.884765322e-14
+ bgidl = 1.758248979e+09 wbgidl = 5.304754484e+1
+ cgidl = 1.546114315e+03 wcgidl = -1.660076109e-3
+ egidl = 4.898457770e-01 wegidl = 6.190923707e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -7.715522461e-01 wkt1 = 7.083407459e-8
+ kt2 = -0.019032
+ at = 5.588748834e+05 wat = -3.346051902e-1
+ ute = -1.515569387e+00 wute = -6.240887629e-8
+ ua1 = 2.2096e-11
+ ub1 = -3.569388362e-18 wub1 = -2.836483427e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.50 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.691765406e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -8.455433763e-08 wvth0 = 9.333710679e-08 pvth0 = 1.301964309e-13
+ k1 = 6.273580940e-01 lk1 = -1.414391571e-07 wk1 = -7.078148731e-08 pk1 = 2.177874483e-13
+ k2 = 1.250383454e-01 lk2 = 3.666195699e-08 wk2 = -3.244789851e-07 pk2 = -5.645193472e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.675729173e+05 lvsat = -1.160728558e+00 wvsat = -2.882850991e-01 pvsat = 1.787285191e-6
+ ua = 2.219459442e-09 lua = 4.027744945e-15 wua = 7.088654414e-16 pua = -6.201905556e-21
+ ub = 3.535876962e-19 lub = -3.961378447e-24 wub = -8.428191912e-25 pub = 6.099714687e-30
+ uc = -8.003679943e-11 luc = 1.835308319e-16 wuc = 8.682878761e-17 puc = -2.826000409e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.899603662e-02 lu0 = 1.057933979e-08 wu0 = 3.499392383e-10 pu0 = -1.629002510e-14
+ a0 = 8.682062231e-01 la0 = -3.004854024e-07 wa0 = 1.422817342e-07 pa0 = 4.626862207e-13
+ keta = -2.223487761e-04 lketa = -4.696243750e-08 wketa = -1.447154362e-08 pketa = 7.231257342e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 7.807165800e-02 lags = 3.160585492e-07 wags = 8.788275113e-08 pags = -4.866656899e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.039819539e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 2.486098478e-08 wvoff = -1.326673700e-08 pvoff = -3.828084492e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.554602573e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -3.935563868e-06 wnfactor = 1.569012509e-07 pnfactor = 6.059965502e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 2.067117695e-02 ltvoff = -9.150727018e-08 wtvoff = -2.741033504e-08 ptvoff = 1.409025286e-13
+ cit = 1.513265333e-05 wcit = -1.560221907e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.164716022e+00 lpclm = 1.157543967e-05 wpclm = 4.629255416e-06 ppclm = -1.782381570e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 7.875866387e-03 lpdiblc2 = -2.551759790e-08 wpdiblc2 = -1.014089072e-08 ppdiblc2 = 3.929189518e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 9.109505333e+08 lpscbe1 = -3.612693517e+03 wpscbe1 = -1.066517809e+03 ppscbe1 = 5.562811026e-3
+ pscbe2 = -4.587929877e-08 lpscbe2 = 4.795353491e-13 wpscbe2 = 9.371885477e-14 ppscbe2 = -7.383866124e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.372007230e-04 lalpha0 = -4.347375954e-10 walpha0 = -1.802329231e-10 palpha0 = 6.694072105e-16
+ alpha1 = 0.0
+ beta0 = 4.083995260e+01 lbeta0 = -1.382760211e-05 wbeta0 = -5.190188217e-06 pbeta0 = 2.129168641e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.703607254e-08 lagidl = -1.514140957e-13 wagidl = 9.240204099e-15 pagidl = 2.331468189e-19
+ bgidl = 1.589234771e+09 lbgidl = 1.330919281e+03 wbgidl = 3.132949461e+02 pbgidl = -2.049344186e-3
+ cgidl = 2.213533951e+03 lcgidl = -5.255662668e-03 wcgidl = -2.687766196e-03 pcgidl = 8.092648353e-9
+ egidl = 1.525886520e+00 legidl = -8.158406432e-06 wegidl = -9.761990207e-07 pegidl = 1.256228159e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -3.783046704e-01 lkt1 = -3.096667360e-06 wkt1 = -5.346869695e-07 pkt1 = 4.768236014e-12
+ kt2 = -0.019032
+ at = 9.890464690e+05 lat = -3.387429168e+00 wat = -9.969816770e-01 pat = 5.215949883e-6
+ ute = -1.476309408e+00 lute = -3.091566275e-07 wute = -1.228612343e-07 pute = 4.760381384e-13
+ ua1 = 2.2096e-11
+ ub1 = -3.390951760e-18 lub1 = -1.405116872e-24 wub1 = -5.584043099e-25 pub1 = 2.163593339e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.51 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.093063217e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 7.093251229e-08 wvth0 = 2.058388430e-07 pvth0 = -3.057027963e-13
+ k1 = 6.237526700e-01 lk1 = -1.274695812e-07 wk1 = -6.522986983e-08 pk1 = 1.962771513e-13
+ k2 = 2.368912380e-01 lk2 = -3.967232609e-07 wk2 = -6.516861804e-07 pk2 = 1.211345064e-12
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.653516055e+04 lvsat = 8.316433416e-02 wvsat = 2.060475545e-01 pvsat = -1.280561091e-7
+ ua = 3.958538769e-09 lua = -2.710491815e-15 wua = -1.968496242e-15 pua = 4.171800023e-21
+ ub = -2.572192094e-18 lub = 7.374847929e-24 wub = 3.568920933e-24 pub = -1.099401360e-29
+ uc = -9.848498936e-11 luc = 2.550101886e-16 wuc = 1.338993559e-16 puc = -4.649796648e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.058214501e-02 lu0 = 4.433804234e-09 wu0 = -2.242139112e-09 pu0 = -6.246758319e-15
+ a0 = 6.025116645e-01 la0 = 7.289747343e-07 wa0 = 6.896066010e-07 pa0 = -1.657978708e-12
+ keta = -6.498185991e-04 lketa = -4.530616293e-08 wketa = -1.381332730e-08 pketa = 6.976224845e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 8.773764353e-02 lags = 2.786067217e-07 wags = 9.665101263e-08 pags = -5.206391959e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-2.924505216e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -2.120829840e-07 wvoff = -1.074301023e-07 pvoff = 3.265645304e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '1.870094371e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 6.465831608e-06 wnfactor = 5.877639136e-06 pnfactor = -1.610560551e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -5.707363990e-03 ltvoff = 1.069902454e-08 wtvoff = 1.734922223e-08 ptvoff = -3.252285199e-14
+ cit = 1.513265333e-05 wcit = -1.560221907e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -4.118600697e-02 leta0 = 4.695473026e-07 weta0 = 1.866017288e-07 peta0 = -7.230070584e-13
+ etab = -1.742655532e-01 letab = 4.039873125e-07 wetab = 1.605476818e-07 petab = -6.220580478e-13
+ dsub = 1.066872821e+00 ldsub = -1.963929431e-06 wdsub = -7.804807418e-07 pdsub = 3.024050682e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.253375859e+00 lpclm = -1.668299137e-06 wpclm = -6.339087899e-07 ppclm = 2.568840339e-12
+ pdiblc1 = 7.711611432e-01 lpdiblc1 = -1.476846965e-06 wpdiblc1 = -5.869104036e-07 ppdiblc1 = 2.274043050e-12
+ pdiblc2 = -3.531850657e-03 lpdiblc2 = 1.868274255e-08 wpdiblc2 = 7.424666354e-09 ppdiblc2 = -2.876761225e-14
+ pdiblcb = 3.548934388e-01 lpdiblcb = -1.471935118e-06 wpdiblcb = -5.849583974e-07 ppdiblcb = 2.266479807e-12
+ drout = -2.757655653e-01 ldrout = 3.238257259e-06 wdrout = 1.286908474e-06 pdrout = -4.986255575e-12
+ pscbe1 = -5.311692445e+08 lpscbe1 = 1.974943774e+03 wpscbe1 = 1.154052457e+03 ppscbe1 = -3.041010524e-3
+ pscbe2 = 1.376797145e-07 lpscbe2 = -2.316824036e-13 wpscbe2 = -1.889245796e-13 ppscbe2 = 3.567436383e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.781846170e-05 lalpha0 = -1.659090859e-10 walpha0 = -7.339839475e-11 palpha0 = 2.554661468e-16
+ alpha1 = -1.899467194e-10 lalpha1 = 7.359675589e-16 walpha1 = 2.924791987e-16 palpha1 = -1.133239903e-21
+ beta0 = 1.025587245e+02 lbeta0 = -2.529631558e-04 wbeta0 = -1.002245063e-04 pbeta0 = 3.895116554e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.786330482e-08 lagidl = 1.000450319e-13 wagidl = 1.132232107e-13 pagidl = -1.697457386e-19
+ bgidl = 2.966981483e+09 lbgidl = -4.007298129e+03 wbgidl = -1.531194103e+03 pbgidl = 5.097313085e-3
+ cgidl = 1.925053268e+03 lcgidl = -4.137915414e-03 wcgidl = -3.300024373e-03 pcgidl = 1.046490389e-8
+ egidl = -4.063873926e+00 legidl = 1.349967939e-05 wegidl = 7.630891755e-06 pegidl = -2.078675233e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -2.028425470e+00 lkt1 = 3.296890689e-06 wkt1 = 2.219489336e-06 pkt1 = -5.903095499e-12
+ kt2 = -0.019032
+ at = 1.766413762e+05 lat = -2.396843955e-01 wat = 3.262200023e-01 pat = 8.907265641e-8
+ ute = -1.617248302e+00 lute = 2.369252119e-07 wute = -1.169916795e-07 pute = 4.532959614e-13
+ ua1 = -4.749579392e-10 lua1 = 1.925885193e-15 wua1 = -4.930380658e-32 pua1 = -3.291384182e-37
+ ub1 = -3.534626259e-18 lub1 = -8.484356564e-25 wub1 = 3.834402295e-25 pub1 = -1.485677513e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.52 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.947797008e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 4.370090871e-08 wvth0 = 8.263529977e-08 pvth0 = -7.474543417e-14
+ k1 = 5.368782874e-01 lk1 = 3.538513637e-08 wk1 = 6.853895696e-08 pk1 = -5.448589143e-14
+ k2 = 1.576593730e-02 lk2 = 1.779822786e-08 wk2 = 8.385982139e-09 pk2 = -2.602621181e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.205052938e+05 lvsat = -2.429600776e-01 wvsat = -2.142979331e-02 pvsat = 2.983729272e-7
+ ua = 4.191991475e-09 lua = -3.148122257e-15 wua = -2.329560282e-15 pua = 4.848650672e-21
+ ub = 1.323788175e-18 lub = 7.144331595e-26 wub = -2.194416571e-24 pub = -1.900611143e-31
+ uc = 7.011423265e-11 luc = -6.104591295e-17 wuc = -2.115764567e-16 puc = 1.826492936e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.063564392e-02 lu0 = -1.441248483e-08 wu0 = -1.707458712e-08 pu0 = 2.155814872e-14
+ a0 = 1.166022590e+00 la0 = -3.273828462e-07 wa0 = -4.900566699e-07 pa0 = 5.534180595e-13
+ keta = 9.491115474e-02 lketa = -2.244447635e-07 wketa = -1.609577318e-07 pketa = 3.455991491e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -7.227527033e-01 lags = 1.797951926e-06 wags = 1.367532876e-06 pags = -2.903034336e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-2.179863479e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.417314491e-07 wvoff = 1.831929900e-07 pvoff = -2.182375184e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '6.890118537e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.944705693e-06 wnfactor = -4.500890962e-06 pnfactor = 3.349987015e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -2.012741666e-03 ltvoff = 3.773085526e-09 wtvoff = 3.099211566e-09 ptvoff = -5.809782001e-15
+ cit = 2.399467194e-05 lcit = -1.661274008e-11 wcit = -2.924791987e-11 pcit = 2.558023072e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 4.486116462e-01 leta0 = -4.486273780e-07 weta0 = -5.675867384e-07 peta0 = 6.907946422e-13
+ etab = 1.446284594e-02 letab = 5.019705542e-08 wetab = -1.300555523e-07 petab = -7.729322514e-14
+ dsub = 8.870340071e-03 ldsub = 1.940201914e-08 wdsub = 8.486272458e-07 pdsub = -2.987515146e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.954494099e-01 lpclm = 1.984968712e-06 wpclm = 2.366887581e-06 ppclm = -3.056452537e-12
+ pdiblc1 = -3.892069132e-01 lpdiblc1 = 6.983789931e-07 wpdiblc1 = 1.199819688e-06 ppdiblc1 = -1.075361180e-12
+ pdiblc2 = 1.055053475e-02 lpdiblc2 = -7.716097123e-09 wpdiblc2 = -1.425933436e-08 ppdiblc2 = 1.188121549e-14
+ pdiblcb = -7.847868775e-01 lpdiblcb = 6.645096031e-07 wpdiblcb = 1.169916795e-06 ppdiblcb = -1.023209229e-12
+ drout = 2.496169776e+00 ldrout = -1.958012731e-06 wdrout = -2.981306476e-06 pdrout = 3.014940172e-12
+ pscbe1 = 6.444177054e+08 lpscbe1 = -2.288115219e+02 wpscbe1 = -6.561116263e+02 ppscbe1 = 3.523230663e-4
+ pscbe2 = 1.406915203e-08 lpscbe2 = 3.795678853e-17 wpscbe2 = 1.410470031e-15 ppscbe2 = -5.844571115e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.408773865e-04 lalpha0 = 2.253121513e-10 walpha0 = 2.479506376e-10 palpha0 = -3.469347492e-16
+ alpha1 = 3.798934388e-10 lalpha1 = -3.322548016e-16 walpha1 = -5.849583974e-16 palpha1 = 5.116046144e-22
+ beta0 = -1.159577660e+02 lbeta0 = 1.566678574e-04 wbeta0 = 2.362463117e-04 pbeta0 = -2.412365401e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.155830798e-08 lagidl = -1.134672351e-14 wagidl = 2.757573301e-14 pagidl = -9.190976898e-21
+ bgidl = 2.042334904e+08 lbgidl = 1.171749257e+03 wbgidl = 2.174264214e+03 pbgidl = -1.848939076e-3
+ cgidl = -1.642687038e+03 lcgidl = 2.550170563e-03 wcgidl = 5.217502413e-03 pcgidl = -5.502051826e-9
+ egidl = 5.301633254e+00 legidl = -4.056900369e-06 wegidl = -6.790078740e-06 pegidl = 6.246798960e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 6.379400959e-03 lkt1 = -5.175545216e-07 wkt1 = -1.451326138e-06 pkt1 = 9.782151890e-13
+ kt2 = -0.019032
+ at = 4.725345396e+04 lat = 2.866203588e-03 wat = 7.551874758e-01 pat = -7.150697696e-7
+ ute = -1.454306515e+00 lute = -6.852546243e-08 wute = 4.294354777e-08 pute = 1.534813843e-13
+ ua1 = 5.524e-10
+ ub1 = -4.333844902e-18 lub1 = 6.497796111e-25 wub1 = -7.668804591e-25 pub1 = 6.707136495e-31
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.53 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-5.746453784e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.362885696e-07 wvth0 = -6.570665711e-07 pvth0 = 5.721978221e-13
+ k1 = 5.829147102e-01 lk1 = -4.878318975e-09 wk1 = 2.066048970e-08 pk1 = -1.261138397e-14
+ k2 = 5.184739692e-02 lk2 = -1.375861672e-08 wk2 = -1.100758034e-07 pk2 = 7.758046580e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.621577801e+05 lvsat = 3.540970468e-01 wvsat = 1.446071540e+00 pvsat = -9.851037387e-7
+ ua = -8.694190006e-09 lua = 8.122132066e-15 wua = 2.430552824e-14 pua = -1.844639775e-20
+ ub = 1.013624510e-17 lub = -7.635931513e-24 wub = -1.981534629e-23 pub = 1.522120402e-29
+ uc = 1.169114993e-11 luc = -9.949084803e-18 wuc = -1.803882766e-17 puc = 1.338128319e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.119653320e-02 lu0 = 2.217393728e-08 wu0 = 6.852001337e-08 pu0 = -5.330288887e-14
+ a0 = 4.524751470e-01 la0 = 2.966857472e-07 wa0 = 1.124022187e-06 pa0 = -8.582553089e-13
+ keta = -4.853074625e-01 lketa = 2.830144391e-07 wketa = 1.018096612e-06 pketa = -6.856017802e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 3.447432368e+00 lags = -1.849291937e-06 wags = -8.688788625e-06 pags = 5.892224448e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-3.634393723e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.713300331e-08 wvoff = -1.764776438e-07 pvoff = 9.633041790e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.063935556e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.347526058e-06 wnfactor = -2.489347783e-06 pnfactor = 1.590691351e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 1.635848925e-02 ltvoff = -1.229439303e-08 wtvoff = -3.158949152e-08 ptvoff = 2.452895772e-14
+ cit = -1.186500000e-05 lcit = 1.475012900e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -2.625933793e-01 leta0 = 1.733925373e-07 weta0 = 9.075794025e-07 peta0 = -5.993856646e-13
+ etab = 3.036900783e-01 letab = -2.027610820e-07 wetab = -9.177019860e-07 petab = 6.115823457e-13
+ dsub = -8.244807420e-01 ldsub = 7.482508756e-07 wdsub = 3.662899848e-06 pdsub = -2.491237969e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.229273684e+00 lpclm = -2.322194106e-06 wpclm = -6.831391685e-06 ppclm = 4.988362509e-12
+ pdiblc1 = 2.388003121e-01 lpdiblc1 = 1.491238739e-07 wpdiblc1 = -1.002779198e-07 ppdiblc1 = 6.170418783e-14
+ pdiblc2 = -4.757742776e-02 lpdiblc2 = 4.312261889e-08 wpdiblc2 = 4.764855928e-08 ppdiblc2 = -4.226342830e-14
+ pdiblcb = -0.025
+ drout = 6.501392062e-02 ldrout = 1.682761797e-07 wdrout = 8.343788724e-07 pdrout = -3.222582343e-13
+ pscbe1 = 2.171666831e+08 lpscbe1 = 1.448622222e+02 wpscbe1 = -7.804351920e+02 ppscbe1 = 4.610564568e-4
+ pscbe2 = 1.609981870e-08 lpscbe2 = -1.738064280e-15 wpscbe2 = 6.078431239e-15 ppscbe2 = -4.141044584e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.050363541e-04 lalpha0 = -3.396040064e-10 walpha0 = -8.105327189e-10 palpha0 = 5.788147943e-16
+ alpha1 = 0.0
+ beta0 = 1.305757067e+02 lbeta0 = -5.895031787e-05 wbeta0 = -1.951898183e-04 pbeta0 = 1.360974991e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.900970465e-08 lagidl = 2.413406034e-14 wagidl = 4.437699541e-15 pagidl = 1.104554717e-20
+ bgidl = 5.910879165e+08 lbgidl = 8.334063764e+02 wbgidl = 4.601843311e+02 pbgidl = -3.498048109e-4
+ cgidl = 3.778797521e+03 lcgidl = -2.191459832e-03 wcgidl = -4.588868505e-03 pcgidl = 3.074600180e-9
+ egidl = 1.727451242e-01 legidl = 4.288251899e-07 wegidl = 4.897698166e-06 pegidl = -3.975330722e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -7.496192309e-01 lkt1 = 1.436418819e-07 wkt1 = -5.777352503e-07 pkt1 = 2.141725982e-13
+ kt2 = -0.019032
+ at = 1.193329324e+05 lat = -6.017450827e-02 wat = -2.202877311e-01 pat = 1.380808464e-7
+ ute = -1.710944302e+00 lute = 1.559299464e-07 wute = 9.551990560e-07 pute = -6.443772832e-13
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.54 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.782713051e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 3.599748048e-08 wvth0 = 3.164037694e-07 pvth0 = -8.450526960e-14
+ k1 = 6.984311726e-01 lk1 = -8.280572453e-08 wk1 = -3.711626561e-07 pk1 = 2.517125102e-13
+ k2 = -1.926915733e-02 lk2 = 3.421661077e-08 wk2 = 1.009238558e-07 pk2 = -6.475990427e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.053382220e+04 lvsat = 2.172729190e-02 wvsat = -6.237696663e-03 pvsat = -5.375927832e-9
+ ua = 2.929858603e-09 lua = 2.805488745e-16 wua = -1.774151785e-15 pua = -8.530456047e-22
+ ub = -5.888109523e-19 lub = -4.008086983e-25 wub = 1.808433741e-24 pub = 6.338020102e-31
+ uc = -5.161753247e-12 luc = 1.419883677e-18 wuc = 8.195147896e-18 puc = -4.316156722e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.660872708e-02 lu0 = -3.329491299e-09 wu0 = -1.369219136e-08 pu0 = 2.157464440e-15
+ a0 = 1.004324241e+00 la0 = -7.559165168e-08 wa0 = -4.888424871e-07 pa0 = 2.297832004e-13
+ keta = -1.403773132e-01 lketa = 5.032456034e-08 wketa = 6.866828687e-08 pketa = -4.511743187e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 6.731453947e-01 lags = 2.224205472e-08 wags = 1.458330132e-07 pags = -6.761130898e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-5.285627237e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.993782023e-09 wvoff = -6.068970537e-08 pvoff = 1.821987462e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.926972956e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.255131088e-06 wnfactor = -2.295057093e-06 pnfactor = 1.459622851e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -6.294780923e-03 ltvoff = 2.987503026e-09 wtvoff = 1.609343369e-08 ptvoff = -7.637943629e-15
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 2.362183104e-02 leta0 = -1.968824363e-08 weta0 = -6.625480182e-08 peta0 = 5.756288963e-14
+ etab = 1.054122412e-02 letab = -5.002864968e-09 wetab = -3.749707003e-08 petab = 1.779610944e-14
+ dsub = 3.008237876e-01 ldsub = -1.087956016e-08 wdsub = -7.901022075e-08 pdsub = 3.305456314e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.582954275e-01 lpclm = 8.678782580e-08 wpclm = 9.542121668e-07 ppclm = -2.638058502e-13
+ pdiblc1 = 3.244687141e-01 lpdiblc1 = 9.133196985e-08 wpdiblc1 = 4.027383038e-07 ppdiblc1 = -2.776305566e-13
+ pdiblc2 = 1.937717598e-02 lpdiblc2 = -2.044956796e-09 wpdiblc2 = -2.421577482e-08 ppdiblc2 = 6.216251490e-15
+ pdiblcb = -0.025
+ drout = 5.487704464e-01 ldrout = -1.580659725e-07 wdrout = -3.555804300e-07 pdrout = 4.804883111e-13
+ pscbe1 = 3.578529221e+08 lpscbe1 = 4.995528530e+01 wpscbe1 = 1.281185187e+02 ppscbe1 = -1.518538764e-4
+ pscbe2 = 1.627824006e-08 lpscbe2 = -1.858427330e-15 wpscbe2 = -8.434294149e-15 ppscbe2 = 5.649239963e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.200845087e-06 lalpha0 = 4.602008251e-12 walpha0 = 6.821611094e-11 palpha0 = -1.398916627e-17
+ alpha1 = 0.0
+ beta0 = 4.496220912e+01 lbeta0 = -1.195452392e-06 wbeta0 = 1.168865031e-06 pbeta0 = 3.633931399e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.953505921e-07 lagidl = -1.879333959e-13 wagidl = -9.061433299e-13 pagidl = 6.253235096e-19
+ bgidl = 1.242353570e+09 lbgidl = 3.940625668e+02 wbgidl = 1.717321899e+03 pbgidl = -1.197869814e-3
+ cgidl = 1.641061823e+03 lcgidl = -7.493433297e-04 wcgidl = -3.407799244e-03 pcgidl = 2.277850856e-9
+ egidl = 3.368809458e+00 legidl = -1.727239809e-06 wegidl = -8.778239257e-06 pegidl = 5.250456664e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.024027736e+00 lkt1 = 3.287578595e-07 wkt1 = 2.188740608e-07 pkt1 = -3.232200431e-13
+ kt2 = -0.019032
+ at = 3.943578152e+04 lat = -6.275890273e-03 wat = 6.612220443e-03 pat = -1.498586090e-8
+ ute = -1.250377861e+00 lute = -1.547681752e-07 wute = -8.596988092e-07 pute = 5.799528167e-13
+ ua1 = 5.533492000e-10 lua1 = -6.403303200e-19
+ ub1 = -8.006595839e-19 lub1 = -1.882296185e-24 wub1 = -1.058592091e-23 pub1 = 7.141262246e-30
+ uc1 = -4.347856431e-10 luc1 = 2.196400749e-16 wuc1 = 5.013354710e-16 puc1 = -3.382009087e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.55 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-5.966792588e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.451061047e-07 wvth0 = -2.942683988e-08 pvth0 = 7.962593756e-14
+ k1 = 4.402571515e-01 lk1 = 3.972366588e-08 wk1 = 5.000616060e-07 pk1 = -1.617705246e-13
+ k2 = 6.573817029e-02 lk2 = -6.127866915e-09 wk2 = -1.682871260e-07 pk2 = 6.300762771e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.664854254e+05 lvsat = 1.152326268e-01 wvsat = 3.075743095e-01 pvsat = -1.543111059e-7
+ ua = 3.861666706e-09 lua = -1.616872514e-16 wua = -7.466718810e-15 pua = 1.848646705e-21
+ ub = -6.158105997e-18 lub = 2.242378730e-24 wub = 1.354432850e-23 pub = -4.936053644e-30
+ uc = 2.488791857e-10 luc = -1.191479459e-16 wuc = -3.821810043e-16 puc = 1.809563651e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 9.059169965e-03 lu0 = 4.999528507e-09 wu0 = 2.140741785e-09 pu0 = -5.356845629e-15
+ a0 = 1.185250763e-01 la0 = 3.448086320e-07 wa0 = 1.267219285e-06 pa0 = -6.036437167e-13
+ keta = -3.411617842e-01 lketa = 1.456168703e-07 wketa = 4.266062779e-07 pketa = -2.149948024e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 5.229230937e+00 lags = -2.140076144e-06 wags = -7.655833886e-06 pags = 3.635059802e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '2.508125825e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.501150206e-07 wvoff = -4.418483999e-07 pvoff = 1.991177910e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.889675575e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.882297507e-07 wnfactor = 2.405102478e-06 pnfactor = -7.710728811e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -9.484175722e-01 leta0 = 4.416416572e-07 weta0 = 1.249024733e-06 peta0 = -5.666687777e-13
+ etab = 6.098984177e-02 letab = -2.894577890e-08 wetab = -1.336073563e-08 petab = 6.341005130e-15
+ dsub = 1.457123012e-01 ldsub = 6.273635131e-08 wdsub = 1.837359667e-07 pdsub = -9.164477743e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.374095369e+00 lpclm = -1.202130827e-06 wpclm = -3.127650509e-06 ppclm = 1.673446176e-12
+ pdiblc1 = 1.735005829e+00 lpdiblc1 = -5.781089451e-07 wpdiblc1 = -8.375439141e-07 ppdiblc1 = 3.110073840e-13
+ pdiblc2 = 5.738295012e-02 lpdiblc2 = -2.008249720e-08 wpdiblc2 = -5.340423413e-08 ppdiblc2 = 2.006909428e-14
+ pdiblcb = 1.493276775e+00 lpdiblcb = -7.205741576e-07 wpdiblcb = -2.337836506e-06 ppdiblcb = 1.109537206e-12
+ drout = -2.722195187e+00 ldrout = 1.394334317e-06 wdrout = 3.117298390e-06 pdrout = -1.167739977e-12
+ pscbe1 = 7.132594476e+08 lpscbe1 = -1.187206517e+02 wpscbe1 = -5.918049225e+02 ppscbe1 = 1.898217887e-4
+ pscbe2 = 4.991142386e-09 lpscbe2 = 3.498429225e-15 wpscbe2 = 1.403897328e-14 ppscbe2 = -5.016572759e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.128203410e-05 lalpha0 = -4.118876621e-11 walpha0 = -2.875816374e-11 palpha0 = 3.203482449e-17
+ alpha1 = -7.591383877e-10 lalpha1 = 3.602870788e-16 walpha1 = 1.168918253e-15 palpha1 = -5.547686028e-22
+ beta0 = 3.554095323e+02 lbeta0 = -1.485337520e-04 wbeta0 = -4.603222410e-04 pbeta0 = 2.226576103e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.179067912e-06 lagidl = 5.118256262e-13 wagidl = 2.753735025e-12 pagidl = -1.111654757e-18
+ bgidl = 7.062135380e+09 lbgidl = -2.368005881e+03 wbgidl = -9.287136651e+03 pbgidl = 4.024846213e-3
+ cgidl = -3.615633147e+03 lcgidl = 1.745484103e-03 wcgidl = 9.742703723e-03 pcgidl = -3.963377852e-9
+ egidl = -1.399748506e+01 legidl = 6.514803569e-06 wegidl = 2.671520617e-05 pegidl = -1.159473253e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 4.237880494e-01 lkt1 = -3.583755123e-07 wkt1 = -1.791363016e-06 pkt1 = 6.308384736e-13
+ kt2 = -0.019032
+ at = 6.985325947e+03 lat = 9.125095941e-03 wat = 3.348236213e-02 pat = -2.773843014e-8
+ ute = -2.820159120e+00 lute = 5.902500105e-07 wute = 2.037343383e-06 pute = -7.949834078e-13
+ ua1 = 5.52e-10
+ ub1 = -8.959456466e-18 lub1 = 1.989868816e-24 wub1 = 1.259198184e-23 pub1 = -3.858970401e-30
+ uc1 = 2.800423226e-11 wuc1 = -2.112665280e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.56 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.196858172e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = 1.713148882e-8
+ k1 = 5.741946117e-01 wk1 = 1.107943015e-8
+ k2 = -3.133503406e-01 wk2 = 3.505501600e-7
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.887126408e+05 wvsat = -3.208359609e-1
+ ua = 3.571354814e-09 wua = -1.372777644e-15
+ ub = -8.942597693e-19 wub = 1.078611345e-24
+ uc = 2.098433423e-11 wuc = -6.872314993e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.150773181e-02 wu0 = -3.517558966e-9
+ a0 = 1.070168137e+00 wa0 = -1.686984135e-7
+ keta = -1.261281697e-02 wketa = 4.607249741e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.729228933e-01 wags = -5.816880151e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-8.099229642e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' wvoff = -2.774990261e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.565351483e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = 1.403501224e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -6.684369526e-03 wtvoff = 1.471162600e-8
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.418357770e+00 wpclm = -2.427743276e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -3.177102117e-03 wpdiblc2 = 6.878425971e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.049994136e+08 wpscbe1 = 2.050290178e+1
+ pscbe2 = 1.495696373e-08 wpscbe2 = 4.342111933e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -7.154207967e-05 walpha0 = 1.411884094e-10
+ alpha1 = 0.0
+ beta0 = 3.420382873e+01 wbeta0 = 5.028088767e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.497105671e-07 wagidl = 4.353735728e-13
+ bgidl = 2.358972902e+09 wbgidl = -8.719447488e+2
+ cgidl = -1.470179744e+03 wcgidl = 2.984401417e-3
+ egidl = -4.141352049e-01 wegidl = 2.011038671e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -5.357664341e-01 wkt1 = -2.922279757e-7
+ kt2 = -0.019032
+ at = 7.376906842e+05 wat = -6.099450450e-1
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -5.161275825e-18 wub1 = 2.167533604e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.57 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.196858172e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = 1.713148882e-8
+ k1 = 5.741946117e-01 wk1 = 1.107943015e-8
+ k2 = -3.133503406e-01 wk2 = 3.505501600e-7
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.887126408e+05 wvsat = -3.208359609e-1
+ ua = 3.571354814e-09 wua = -1.372777644e-15
+ ub = -8.942597693e-19 wub = 1.078611345e-24
+ uc = 2.098433423e-11 wuc = -6.872314993e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.150773181e-02 wu0 = -3.517558966e-9
+ a0 = 1.070168137e+00 wa0 = -1.686984135e-7
+ keta = -1.261281697e-02 wketa = 4.607249741e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.729228933e-01 wags = -5.816880151e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-8.099229642e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' wvoff = -2.774990261e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.565351483e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = 1.403501224e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -6.684369526e-03 wtvoff = 1.471162600e-8
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.418357770e+00 wpclm = -2.427743276e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -3.177102117e-03 wpdiblc2 = 6.878425971e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.049994136e+08 wpscbe1 = 2.050290178e+1
+ pscbe2 = 1.495696373e-08 wpscbe2 = 4.342111933e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -7.154207967e-05 walpha0 = 1.411884094e-10
+ alpha1 = 0.0
+ beta0 = 3.420382873e+01 wbeta0 = 5.028088767e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.497105671e-07 wagidl = 4.353735728e-13
+ bgidl = 2.358972902e+09 wbgidl = -8.719447488e+2
+ cgidl = -1.470179744e+03 wcgidl = 2.984401417e-3
+ egidl = -4.141352049e-01 wegidl = 2.011038671e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -5.357664341e-01 wkt1 = -2.922279757e-7
+ kt2 = -0.019032
+ at = 7.376906842e+05 wat = -6.099450450e-1
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -5.161275825e-18 wub1 = 2.167533604e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.58 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.504859441e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 2.425386795e-07 wvth0 = 6.455740107e-08 pvth0 = -3.734600886e-13
+ k1 = 6.149861467e-01 lk1 = -3.212170216e-07 wk1 = -5.173121229e-08 pk1 = 4.946086850e-13
+ k2 = -3.253686025e-01 lk2 = 9.463900518e-08 wk2 = 3.690558316e-07 pk2 = -1.457247616e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.694375778e+05 lvsat = -6.356765889e-01 wvsat = -4.451358960e-01 pvsat = 9.788122688e-7
+ ua = 2.999199827e-09 lua = 4.505491656e-15 wua = -4.917756849e-16 pua = -6.937538030e-21
+ ub = -6.297090387e-19 lub = -2.083231183e-24 wub = 6.712571881e-25 pub = 3.207751042e-30
+ uc = 5.161629932e-11 luc = -2.412144723e-16 wuc = -1.158901272e-16 puc = 3.714210796e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.008677632e-02 lu0 = 1.118945615e-08 wu0 = -1.329577377e-09 pu0 = -1.722947982e-14
+ a0 = 9.951455548e-01 la0 = 5.907728286e-07 wa0 = -5.317894100e-08 pa0 = -9.096696384e-13
+ keta = -1.592710401e-02 lketa = 2.609868472e-08 wketa = 9.710575668e-09 pketa = -4.018665034e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.614313840e-01 lags = 9.049103857e-08 wags = -4.047422156e-08 pags = -1.393377392e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-5.962025352e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.682962890e-07 wvoff = -6.065848877e-08 pvoff = 2.591419526e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.868947369e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 1.335850383e-05 wnfactor = 2.752466391e-06 pnfactor = -2.056937077e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -2.172023005e-02 ltvoff = 1.184013873e-07 wtvoff = 3.786378389e-08 ptvoff = -1.823139826e-13
+ cit = 1.507198395e-05 lcit = -7.931284484e-11 wcit = -1.550880060e-11 pcit = 1.221256012e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.090490658e+00 lpclm = -1.316737764e-05 wpclm = -5.002486808e-06 ppclm = 2.027507542e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -7.504160582e-03 lpdiblc2 = 3.407385459e-08 wpdiblc2 = 1.354121329e-08 ppdiblc2 = -5.246678501e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.056864437e+08 lpscbe1 = -5.410087773e+00 wpscbe1 = 1.944501547e+01 ppscbe1 = 8.330431512e-6
+ pscbe2 = 1.497442050e-08 lpscbe2 = -1.374650227e-16 wpscbe2 = 1.654126612e-17 ppscbe2 = 2.116680921e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.009520481e-04 lalpha0 = 1.019051737e-09 walpha0 = 3.404533612e-10 palpha0 = -1.569131789e-15
+ alpha1 = 2.014396791e-10 lalpha1 = -1.586256897e-15 walpha1 = -3.101760121e-16 palpha1 = 2.442512025e-21
+ beta0 = -3.839398009e+01 lbeta0 = 5.716787054e-04 wbeta0 = 1.168139044e-04 pbeta0 = -8.802685838e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.825707221e-07 lagidl = -5.286994237e-13 wagidl = 3.319919080e-13 pagidl = 8.140892579e-19
+ bgidl = 2.262080416e+09 lbgidl = 7.629895674e+02 wbgidl = -7.227500870e+02 pbgidl = -1.174848284e-3
+ cgidl = -3.299252030e+03 lcgidl = 1.440321262e-02 wcgidl = 5.800799607e-03 pcgidl = -2.217800919e-8
+ egidl = 5.529057876e-01 legidl = -7.615061000e-06 wegidl = 5.219928187e-07 pegidl = 1.172564047e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -8.224755293e-01 lkt1 = 2.257719441e-06 wkt1 = 1.492455423e-07 pkt1 = -3.476427365e-12
+ kt2 = -0.019032
+ at = 8.757977281e+05 lat = -1.087537729e+00 wat = -8.226017189e-01 pat = 1.674586244e-6
+ ute = -1.262602388e+00 lute = -2.311176299e-06 wute = -4.519264496e-07 pute = 3.558740020e-12
+ ua1 = 2.2096e-11
+ ub1 = -3.797730637e-18 lub1 = -1.073737294e-23 wub1 = 6.795217850e-26 pub1 = 1.653336390e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.59 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-6.646181862e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -4.776245353e-07 wvth0 = -1.709309693e-07 pvth0 = 5.389631513e-13
+ k1 = 5.094331513e-01 lk1 = 8.775861433e-08 wk1 = 1.107988678e-07 pk1 = -1.351303633e-13
+ k2 = -5.981118917e-01 lk2 = 1.151410153e-06 wk2 = 6.340482987e-07 pk2 = -1.172464575e-12
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.120844454e+05 lvsat = 7.489238581e-01 wvsat = 1.051150279e-01 pvsat = -1.153189961e-6
+ ua = 3.548390458e-09 lua = 2.377597638e-15 wua = -1.336951513e-15 pua = -3.662819765e-21
+ ub = -9.844732780e-19 lub = -7.086616611e-25 wub = 1.124157851e-24 pub = 1.452942134e-30
+ uc = 6.096499929e-11 luc = -2.774369452e-16 wuc = -1.116210988e-16 puc = 3.548803021e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.101884943e-02 lu0 = 7.578045679e-09 wu0 = -2.914574823e-09 pu0 = -1.108824872e-14
+ a0 = 1.553080492e+00 la0 = -1.571001879e-06 wa0 = -7.740754772e-07 pa0 = 1.883516081e-12
+ keta = -2.139603482e-01 lketa = 7.933982925e-07 wketa = 3.146413729e-07 pketa = -1.221671517e-12
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.348510155e+00 lags = -4.508964369e-06 wags = -1.844681458e-06 pags = 6.851243620e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-8.178467558e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -8.241801929e-08 wvoff = -2.652980034e-08 pvoff = 1.269069364e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '9.183185441e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.110664300e-05 wnfactor = -5.383029241e-06 pnfactor = 1.095242061e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 1.712209197e-02 ltvoff = -3.209707361e-08 wtvoff = -1.780348274e-08 ptvoff = 3.337440875e-14
+ cit = -1.135086139e-05 lcit = 2.306511174e-11 wcit = 2.517699097e-11 pcit = -3.551556680e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -7.593611893e-02 leta0 = 6.041901158e-07 weta0 = 2.401098239e-07 peta0 = -9.303295236e-13
+ etab = 6.518102809e-02 letab = -5.237724114e-07 wetab = -2.081512063e-07 petab = 8.065026640e-13
+ dsub = -2.476047448e-02 ldsub = 2.265712934e-06 wdsub = 9.004118396e-07 pdsub = -3.488735714e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.621645791e+00 lpclm = -7.476191322e-06 wpclm = -2.740765358e-06 ppclm = 1.151180949e-11
+ pdiblc1 = 3.917704598e-01 lpdiblc1 = -6.859823528e-09 wpdiblc1 = -2.726146913e-09 ppdiblc1 = 1.056272883e-14
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 7.120380547e-01 ldrout = -5.890866469e-07 wdrout = -2.341075885e-07 pdrout = 9.070732625e-13
+ pscbe1 = 3.696678366e+08 lpscbe1 = -6.407723924e+02 wpscbe1 = -2.330528773e+02 ppscbe1 = 9.866587667e-4
+ pscbe2 = 1.447215109e-08 lpscbe2 = 1.808628007e-15 wpscbe2 = 7.899336841e-16 ppscbe2 = -2.784918171e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.853471021e-04 lalpha0 = -2.415002950e-09 walpha0 = -1.024266525e-09 palpha0 = 3.718611882e-15
+ alpha1 = -4.028793582e-10 lalpha1 = 7.552376448e-16 walpha1 = 6.203520242e-16 palpha1 = -1.162911905e-21
+ beta0 = 2.111793498e+02 lbeta0 = -3.953181187e-04 wbeta0 = -2.674781107e-04 pbeta0 = 6.087092579e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.415234233e-07 lagidl = 8.717871268e-14 wagidl = 5.807978466e-13 pagidl = -1.499342319e-19
+ bgidl = 3.272749501e+09 lbgidl = -3.152948870e+03 wbgidl = -2.002014475e+03 pbgidl = 3.781789514e-3
+ cgidl = -1.016507215e+03 lcgidl = 5.558489565e-03 wcgidl = 1.229378693e-03 pcgidl = -4.465581713e-9
+ egidl = -2.470753358e+00 legidl = 4.100408724e-06 wegidl = 5.177811076e-06 pegidl = -6.313792952e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 4.705040162e-01 lkt1 = -2.752059106e-06 wkt1 = -1.628352291e-06 pkt1 = 3.411053198e-12
+ kt2 = -0.019032
+ at = 3.443156213e+05 lat = 9.717428428e-01 wat = 6.803587046e-02 pat = -1.776278159e-6
+ ute = -2.268527005e+00 lute = 1.586379225e-06 wute = 8.858446624e-07 pute = -1.624587931e-12
+ ua1 = -4.426235773e-11 lua1 = 2.571120929e-16 wua1 = -6.631833336e-16 pua1 = 2.569570144e-21
+ ub1 = -5.909546164e-18 lub1 = -2.554932493e-24 wub1 = 4.040332400e-24 pub1 = 1.141979490e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.60 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.227140619e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 6.201993296e-09 wvth0 = 1.256485172e-07 pvth0 = -1.700475421e-14
+ k1 = 5.613222159e-01 lk1 = -9.512626104e-09 wk1 = 3.090029374e-08 pk1 = 1.464750362e-14
+ k2 = 1.473811222e-02 lk2 = 2.561536001e-09 wk2 = 9.968623091e-09 pk2 = -2.564814635e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.375736987e+05 lvsat = -2.361582961e-01 wvsat = -6.636300549e-01 pvsat = 2.878995712e-7
+ ua = 3.513168799e-09 lua = 2.443624159e-15 wua = -1.284311842e-15 pua = -3.761498093e-21
+ ub = -1.772636327e-19 lub = -2.221856862e-24 wub = 1.168969990e-25 pub = 3.341153327e-30
+ uc = -1.632522026e-10 luc = 1.428806216e-16 wuc = 1.477602469e-16 puc = -1.313559686e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.188165071e-02 lu0 = 5.960638397e-09 wu0 = -3.595223383e-09 pu0 = -9.812304928e-15
+ a0 = 5.026427648e-01 la0 = 3.981486846e-07 wa0 = 5.314129311e-07 pa0 = -5.637524895e-13
+ keta = 2.591947894e-01 lketa = -9.357832834e-08 wketa = -4.139210153e-07 pketa = 1.440915357e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -9.620606373e-01 lags = -1.775683611e-07 wags = 1.736018275e-06 pags = 1.388638994e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.139044748e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -2.220624369e-08 wvoff = 2.292813800e-08 pvoff = 3.419308521e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.185031520e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 1.374963392e-07 wnfactor = 1.204187207e-06 pnfactor = -1.395975345e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.586213028e-06 lcit = 6.634901914e-12 wcit = 1.168122048e-11 pcit = -1.021639543e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 3.182868228e-01 leta0 = -1.348201654e-07 weta0 = -3.669130477e-07 peta0 = 2.075955514e-13
+ etab = -2.144751513e-01 letab = 4.710625170e-10 wetab = 2.224622601e-07 petab = -7.253401795e-16
+ dsub = 1.271023372e+00 ldsub = -1.633634649e-07 wdsub = -1.094830945e-06 pdsub = 2.515464097e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.522520662e+00 lpclm = 2.167063111e-06 wpclm = 5.180204586e-06 ppclm = -3.336840766e-12
+ pdiblc1 = 2.686891478e-01 lpdiblc1 = 2.238684039e-07 wpdiblc1 = 1.867939649e-07 ppdiblc1 = -3.447116728e-13
+ pdiblc2 = 2.604457374e-03 lpdiblc2 = -2.464081793e-09 wpdiblc2 = -2.023996207e-09 ppdiblc2 = 3.794183289e-15
+ pdiblcb = -0.025
+ drout = 1.056200202e+00 ldrout = -1.234253008e-06 wdrout = -7.640470865e-07 pdrout = 1.900497845e-12
+ pscbe1 = 2.991295334e+07 lpscbe1 = -3.867888327e+00 wpscbe1 = 2.901003329e+02 ppscbe1 = 5.955758974e-6
+ pscbe2 = 1.480125856e-08 lpscbe2 = 1.191683154e-15 wpscbe2 = 2.831753268e-16 ppscbe2 = -1.834948954e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.049510260e-03 lalpha0 = 8.371606617e-10 walpha0 = 1.647059902e-09 palpha0 = -1.289056638e-15
+ alpha1 = 0.0
+ beta0 = -9.508645114e+00 lbeta0 = 1.838359660e-05 wbeta0 = 7.233638114e-05 pbeta0 = -2.830698851e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.028809658e-07 lagidl = 5.771195617e-13 wagidl = 9.890848290e-13 pagidl = -9.153090090e-19
+ bgidl = 1.524633757e+09 lbgidl = 1.240689036e+02 wbgidl = 1.411171648e+02 pbgidl = -2.357250583e-4
+ cgidl = 2.756639714e+03 lcgidl = -1.514651668e-03 wcgidl = -1.556563321e-03 pcgidl = 7.569451873e-10
+ egidl = -2.751656863e+00 legidl = 4.626990435e-06 wegidl = 5.610345169e-06 pegidl = -7.124621363e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.100738476e+00 lkt1 = 1.933920699e-07 wkt1 = 2.534095398e-07 pkt1 = -1.164975288e-13
+ kt2 = -0.019032
+ at = 1.644827130e+06 lat = -1.466196031e+00 wat = -1.704750080e+00 pat = 1.546986383e-6
+ ute = -1.557117678e+00 lute = 2.527712995e-07 wute = 2.012517647e-07 pute = -3.412500844e-13
+ ua1 = -3.089911629e-10 lua1 = 7.533727111e-16 wua1 = 1.326366667e-15 pua1 = -1.160040287e-21
+ ub1 = -1.049236659e-17 lub1 = 6.036022682e-24 wub1 = 8.715986607e-24 pub1 = -7.623001886e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.61 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.302991059e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 3.387922552e-07 wvth0 = 4.644371948e-07 pvth0 = -3.133093316e-13
+ k1 = 4.610128395e-01 lk1 = 7.821795450e-08 wk1 = 2.083645026e-07 pk1 = -1.405626935e-13
+ k2 = -3.962219969e-02 lk2 = 5.010506479e-08 wk2 = 3.076871561e-08 pk2 = -2.075657555e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.426811871e+06 lvsat = -9.264260020e-01 wvsat = -1.462556374e+00 pvsat = 9.866405298e-7
+ ua = 2.295241408e-08 lua = -1.455793977e-14 wua = -2.442378615e-14 pua = 1.647628614e-20
+ ub = -1.391389109e-17 lub = 9.792197509e-24 wub = 1.721695721e-23 pub = -1.161455933e-29
+ uc = 6.875872891e-12 luc = -5.913393293e-18 wuc = -1.062428334e-17 puc = 7.167141543e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 7.537561653e-02 lu0 = -4.082518411e-08 wu0 = -6.478343649e-08 pu0 = 4.370290626e-14
+ a0 = 1.503858504e+00 la0 = -4.775146006e-07 wa0 = -4.948936998e-07 pa0 = 3.338552899e-13
+ keta = 8.835203133e-01 lketa = -6.396134316e-07 wketa = -1.089618922e-06 pketa = 7.350569245e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -7.576570838e+00 lags = 5.607482260e-06 wags = 8.285927415e-06 pags = -5.589686634e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-3.271018151e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.642561502e-07 wvoff = 2.712301735e-07 pvoff = -1.829718751e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.560374232e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.065378397e-06 wnfactor = -1.713966070e-06 pnfactor = 1.156241511e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -4.156885200e-03 ltvoff = 3.635611796e-9
+ cit = -1.186500000e-05 lcit = 1.475012900e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 6.947492836e-01 leta0 = -4.640742614e-07 weta0 = -5.665330005e-07 peta0 = 3.821831622e-13
+ etab = -9.217337757e-01 letab = 6.190394554e-07 wetab = 9.692007626e-07 petab = -6.538228345e-13
+ dsub = 3.846828652e+00 ldsub = -2.416162763e-06 wdsub = -3.529963672e-06 pdsub = 2.381313493e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.083660311e+00 lpclm = 3.532435848e-06 wpclm = 5.968830827e-06 ppclm = -4.026573276e-12
+ pdiblc1 = 7.625258158e-01 lpdiblc1 = -2.080411459e-07 wpdiblc1 = -9.067083554e-07 ppdiblc1 = 6.116654566e-13
+ pdiblc2 = -2.320499255e-02 lpdiblc2 = 2.010886311e-08 wpdiblc2 = 1.011998103e-08 ppdiblc2 = -6.826939205e-15
+ pdiblcb = -0.025
+ drout = -3.394491394e+00 ldrout = 2.658321861e-06 wdrout = 6.161311317e-06 pdrout = -4.156420615e-12
+ pscbe1 = -1.132897054e+09 lpscbe1 = 1.013125744e+03 wpscbe1 = 1.298387551e+03 ppscbe1 = -8.758922416e-4
+ pscbe2 = 2.520157653e-08 lpscbe2 = -7.904434946e-15 wpscbe2 = -7.936419066e-15 ppscbe2 = 5.353908302e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.131780585e-04 lalpha0 = 3.680845179e-10 walpha0 = 7.573097608e-10 palpha0 = -5.108811646e-16
+ alpha1 = 0.0
+ beta0 = -1.097040904e+02 lbeta0 = 1.060145330e-04 wbeta0 = 1.747920522e-04 pbeta0 = -1.179147184e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.470608576e-07 lagidl = -7.877955702e-14 wagidl = -2.512770879e-13 pagidl = 1.695115235e-19
+ bgidl = 1.254620138e+09 lbgidl = 3.602228148e+02 wbgidl = -5.615199298e+02 pbgidl = 3.788013447e-4
+ cgidl = 2.761297126e+03 lcgidl = -1.518725041e-03 wcgidl = -3.022125468e-03 pcgidl = 2.038725841e-9
+ egidl = 1.055513705e+01 legidl = -7.011131521e-06 wegidl = -1.108906739e-05 pegidl = 7.480684862e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.466212548e+00 lkt1 = 5.130356937e-07 wkt1 = 5.256722735e-07 pkt1 = -3.546185157e-13
+ kt2 = -0.019032
+ at = -2.056111163e+05 lat = 1.521972591e-01 wat = 2.800598154e-01 pat = -1.889283515e-7
+ ute = -5.540537069e-01 lute = -6.245084494e-07 wute = -8.261764554e-07 pute = 5.573386368e-13
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.62 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.727870920e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.888334114e-8
+ k1 = 4.573845300e-01 lk1 = 8.066561206e-8
+ k2 = 4.627449637e-02 lk2 = -7.840846369e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.648283320e+04 lvsat = 1.823596718e-2
+ ua = 1.777659360e-09 lua = -2.734502297e-16
+ ub = 5.856522500e-19 lub = 1.080557415e-26
+ uc = 1.604763834e-13 luc = -1.383186809e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.771651580e-02 lu0 = -1.928354759e-9
+ a0 = 6.868520000e-01 la0 = 7.363798680e-8
+ keta = -9.578160900e-02 lketa = 2.102364523e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 7.678547025e-01 lags = -2.166720922e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.227039305e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 5.838872834e-9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.436478700e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -3.071984710e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 4.156885200e-03 ltvoff = -1.972857716e-9
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.940646740e-02 leta0 = 1.769520823e-8
+ etab = -1.381074850e-02 letab = 6.554581238e-9
+ dsub = 2.495116523e-01 ldsub = 1.058728554e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.277995808e+00 lpclm = -8.453736934e-8
+ pdiblc1 = 5.860217405e-01 lpdiblc1 = -8.897149673e-8
+ pdiblc2 = 3.650563609e-03 lpdiblc2 = 1.992104925e-9
+ pdiblcb = -0.025
+ drout = 3.178434729e-01 ldrout = 1.539807603e-7
+ pscbe1 = 4.410577874e+08 lpscbe1 = -4.866419185e+1
+ pscbe2 = 1.080070008e-08 lpscbe2 = 1.810396309e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.910119943e-05 lalpha0 = -4.483069431e-12
+ alpha1 = 0.0
+ beta0 = 4.572131294e+01 lbeta0 = 1.164555946e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.931321224e-07 lagidl = 2.181746273e-13 wagidl = 1.009741959e-28 pagidl = -2.407412430e-35
+ bgidl = 2.357645400e+09 lbgidl = -3.838780268e+2
+ cgidl = -5.720880000e+02 lcgidl = 7.299765648e-4
+ egidl = -2.332101090e+00 legidl = 1.682599328e-06 pegidl = -1.009741959e-28
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -8.818828930e-01 lkt1 = 1.188469082e-7
+ kt2 = -0.019032
+ at = 4.373000000e+04 lat = -1.600825800e-2
+ ute = -1.808697800e+00 lute = 2.218744559e-7
+ ua1 = 5.533492000e-10 lua1 = -6.403303200e-19
+ ub1 = -7.675544900e-18 lub1 = 2.755501450e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.63 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-6.717857379e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -6.681858378e-08 wvth0 = 8.622181619e-08 pvth0 = -4.092087396e-14
+ k1 = 5.225080797e-01 lk1 = 4.975797538e-08 wk1 = 3.734119558e-07 pk1 = -1.772213142e-13
+ k2 = 8.659299677e-03 lk2 = 1.001132598e-08 wk2 = -8.039730939e-08 pk2 = 3.815656304e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.146068784e+05 lvsat = -7.104770465e-02 wvsat = -2.792300954e-01 pvsat = 1.325226033e-7
+ ua = -5.023024349e-09 lua = 2.954154258e-15 wua = 6.213892938e-15 pua = -2.949113588e-21
+ ub = 8.268643517e-18 lub = -3.635542081e-24 wub = -8.669922691e-24 pub = 4.114745309e-30
+ uc = -1.708189661e-11 luc = 6.800043412e-18 wuc = 2.734480638e-17 puc = -1.297784511e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 7.651223734e-03 lu0 = 2.848632856e-09 wu0 = 4.308691761e-09 pu0 = -2.044905110e-15
+ a0 = 2.036984989e-01 la0 = 3.029426384e-07 wa0 = 1.136069590e-06 pa0 = -5.391786273e-13
+ keta = 2.445806335e-01 lketa = -1.405122751e-07 wketa = -4.753175539e-07 pketa = 2.255857111e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -5.433737334e+00 lags = 2.921608371e-06 wags = 8.762962005e-06 pags = -4.158901767e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-2.037444327e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 5.874445205e-08 wvoff = 2.580766740e-07 pvoff = -1.224831895e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '-1.005208075e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 1.800826072e-06 wnfactor = 8.402428743e-06 pnfactor = -3.987792681e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.895075816e-05 lcit = 1.848602982e-11 wcit = 5.997622161e-11 pcit = -2.846471478e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 6.194724414e-01 leta0 = -2.855167219e-07 weta0 = -1.165206038e-06 peta0 = 5.530067857e-13
+ etab = 7.583135778e-02 letab = -3.598956240e-08 wetab = -3.621364261e-08 petab = 1.718699478e-14
+ dsub = 3.006359110e-01 ldsub = -1.367628763e-08 wdsub = -5.481478793e-08 pdsub = 2.601509835e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.728204398e+00 lpclm = 1.342205248e-06 wpclm = 4.728850263e-06 ppclm = -2.244312335e-12
+ pdiblc1 = 7.690301627e-01 lpdiblc1 = -1.758272939e-07 wpdiblc1 = 6.498615536e-07 ppdiblc1 = -3.084242933e-13
+ pdiblc2 = 8.637866868e-03 lpdiblc2 = -3.748692020e-10 wpdiblc2 = 2.165325007e-08 ppdiblc2 = -1.027663249e-14
+ pdiblcb = -1.583030326e+00 lpdiblcb = 7.394411929e-07 wpdiblcb = 2.399048864e-06 ppdiblcb = -1.138588591e-12
+ drout = -6.977072743e-01 ldrout = 6.359611450e-7
+ pscbe1 = 3.903948902e+09 lpscbe1 = -1.692152315e+03 wpscbe1 = -5.504815781e+03 ppscbe1 = 2.612585570e-3
+ pscbe2 = -5.650026241e-08 lpscbe2 = 3.375143310e-14 wpscbe2 = 1.087231924e-13 ppscbe2 = -5.160002712e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.793161463e-05 lalpha0 = 3.207670412e-11 walpha0 = 1.702044957e-10 palpha0 = -8.077905367e-17
+ alpha1 = 0.0
+ beta0 = -4.884413343e+00 lbeta0 = 2.518203364e-05 wbeta0 = 9.445693526e-05 pbeta0 = -4.482926148e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.072282781e-06 lagidl = -4.298512858e-13 wagidl = -7.128857667e-13 pagidl = 3.383355849e-19
+ bgidl = 3.828950666e+09 lbgidl = -1.082159506e+03 wbgidl = -4.308691761e+03 pbgidl = 2.044905110e-3
+ cgidl = 1.153605674e+03 lcgidl = -8.903765269e-05 wcgidl = 2.399048864e-03 pcgidl = -1.138588591e-9
+ egidl = -5.967441155e-01 legidl = 8.589989077e-07 wegidl = 6.080798865e-06 pegidl = -2.885947141e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.510350521e-01 lkt1 = -2.280134771e-07 wkt1 = -9.062527038e-07 pkt1 = 4.301075332e-13
+ kt2 = -0.019032
+ at = -2.430606528e+03 lat = 5.899565858e-03 wat = 4.798097729e-02 pat = -2.277177182e-8
+ ute = -8.831696514e-01 lute = -2.173812034e-07 wute = -9.452252526e-07 pute = 4.486039049e-13
+ ua1 = 5.52e-10
+ ub1 = -7.817616000e-19 lub1 = -5.162881046e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.64 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.341384114e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = 3.215923842e-8
+ k1 = 6.285415147e-01 wk1 = -4.543026224e-8
+ k2 = 9.090363253e-03 wk2 = 1.527760591e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.363752817e+05 wvsat = 3.291279606e-1
+ ua = 1.986849924e-09 wua = 2.747842021e-16
+ ub = 5.757518406e-19 wub = -4.499008472e-25
+ uc = -8.450228594e-11 wuc = 4.096141578e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.579932466e-02 wu0 = 2.418019959e-9
+ a0 = 1.006639111e+00 wa0 = -1.026411860e-7
+ keta = -9.711576893e-03 wketa = 1.590551914e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 9.354043521e-02 wags = 2.437276083e-8
+ b0 = -2.962303653e-07 wb0 = 3.080191489e-13
+ b1 = -9.769776520e-10 wb1 = 1.015857455e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.034038269e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' wvoff = -4.446482811e-9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.016343176e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = -3.285892359e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 2.153678513e-02 wtvoff = -1.463261773e-8
+ cit = -1.079592000e-05 wcit = 1.642453443e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.795808282e+00 wpclm = 2.993925728e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.022420423e-02 wpdiblc2 = -7.056198767e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.219288719e+08 wpscbe1 = 2.899718705e+0
+ pscbe2 = 1.501243070e-08 wpscbe2 = -1.425321098e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.072399077e-04 walpha0 = -1.486879859e-10
+ alpha1 = 0.0
+ beta0 = 4.331374970e+01 wbeta0 = -4.444370615e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.376309236e-07 wagidl = -1.753417598e-13
+ bgidl = 9.470081040e+08 wbgidl = 5.962105999e+2
+ cgidl = 2.031836800e+03 wcgidl = -6.569813773e-4
+ egidl = 2.881090477e+00 wegidl = -1.415323812e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.220269389e+00 wkt1 = 4.195154585e-7
+ kt2 = -0.019032
+ at = -4.818525144e+05 wat = 6.581310947e-1
+ ute = -2.016393109e+00 wute = 4.786109334e-7
+ ua1 = 2.2096e-11
+ ub1 = -5.215151650e-18 wub1 = 2.223553471e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.65 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.544341504e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 4.033696945e-07 wvth0 = 5.326266666e-08 pvth0 = -4.194221948e-13
+ k1 = 6.572126149e-01 lk1 = -5.698266471e-07 wk1 = -7.524235749e-08 pk1 = 5.925034683e-13
+ k2 = -5.513545684e-04 lk2 = 1.916252850e-07 wk2 = 2.530302553e-08 pk2 = -1.992512049e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.440883843e+05 lvsat = 4.128214828e+00 wvsat = 5.451072138e-01 pvsat = -4.292501266e-6
+ ua = 1.813433241e-09 lua = 3.446587204e-15 wua = 4.551021752e-16 pua = -3.583747589e-21
+ ub = 8.596848758e-19 lub = -5.643055501e-24 wub = -7.451332814e-25 pub = 5.867626538e-30
+ uc = -1.103530910e-10 luc = 5.137744108e-16 wuc = 6.784097951e-17 puc = -5.342205773e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.427330898e-02 lu0 = 3.032895119e-08 wu0 = 4.004764957e-09 pu0 = -3.153592213e-14
+ a0 = 1.071416103e+00 la0 = -1.287416801e-06 wa0 = -1.699960430e-07 pa0 = 1.338650840e-12
+ keta = -1.071537636e-02 lketa = 1.995011298e-08 wketa = 2.634298590e-09 pketa = -2.074404768e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 7.815875277e-02 lags = 3.057047858e-07 wags = 4.036657270e-08 pags = -3.178706134e-13
+ b0 = -4.906216682e-07 lb0 = 3.863449388e-12 wb0 = 5.101464481e-13 pb0 = -4.017199220e-18
+ b1 = -1.618086670e-09 lb1 = 1.274178529e-14 wb1 = 1.682480047e-15 pb1 = -1.324885738e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.005976456e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.577173158e-08 wvoff = -7.364338939e-09 pvoff = 5.799122341e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.223716288e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -4.121457665e-06 wnfactor = -5.442149689e-07 pnfactor = 4.285475194e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 3.077145003e-02 ltvoff = -1.835352711e-07 wtvoff = -2.423478535e-08 ptvoff = 1.908392408e-13
+ cit = -2.116146597e-05 lcit = 2.060110799e-10 wcit = 2.720258767e-11 pcit = -2.142094969e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.685278872e+00 lpclm = 3.755247219e-05 wpclm = 4.958589690e-06 ppclm = -3.904691037e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 1.467738085e-02 lpdiblc2 = -8.850510400e-08 wpdiblc2 = -1.168659400e-08 ppdiblc2 = 9.202725312e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.200988555e+08 lpscbe1 = 3.637084414e+01 wpscbe1 = 4.802562448e+00 ppscbe1 = -3.781825825e-5
+ pscbe2 = 1.502142592e-08 lpscbe2 = -1.787764152e-16 wpscbe2 = -2.360640558e-17 ppscbe2 = 1.858910014e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.010770973e-04 lalpha0 = -1.864976610e-09 walpha0 = -2.462595204e-10 palpha0 = 1.939195219e-15
+ alpha1 = 0.0
+ beta0 = 4.611859803e+01 lbeta0 = -5.574523855e-05 wbeta0 = -7.360840686e-06 pbeta0 = 5.796367607e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.482893461e-07 lagidl = -2.199291885e-12 wagidl = -2.904039449e-13 pagidl = 2.286814905e-18
+ bgidl = 5.707387853e+08 lbgidl = 7.478202201e+03 wbgidl = 9.874539324e+02 pbgidl = -7.775804736e-3
+ cgidl = 2.446458639e+03 lcgidl = -8.240443197e-03 wcgidl = -1.088103507e-03 pcgidl = 8.568379874e-9
+ egidl = 3.774303256e+00 legidl = -1.775224669e-05 wegidl = -2.344082887e-06 pegidl = 1.845871510e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.485026164e+00 lkt1 = 5.261935003e-06 wkt1 = 6.948084942e-07 pkt1 = -5.471338969e-12
+ kt2 = -0.019032
+ at = -8.971999414e+05 lat = 8.254863972e+00 wat = 1.090007688e+00 pat = -8.583374539e-6
+ ute = -2.318445118e+00 lute = 6.003162869e-06 wute = 7.926834047e-07 pute = -6.242064738e-12
+ ua1 = 2.2096e-11
+ ub1 = -6.618439263e-18 lub1 = 2.788978000e-23 wub1 = 3.682686319e-24 pub1 = -2.899968168e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.66 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.116509405e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -7.209909701e-07 wvth0 = -7.980268039e-08 pvth0 = 6.284141870e-13
+ k1 = 4.609451442e-01 lk1 = 9.757011772e-07 wk1 = 1.084400059e-07 pk1 = -8.539216704e-13
+ k2 = 6.205204052e-02 lk2 = -3.013514100e-07 wk2 = -3.378260332e-08 pk2 = 2.660244881e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.253141520e+05 lvsat = -1.143062384e+00 wvsat = -1.912973343e-01 pvsat = 1.506389989e-6
+ ua = 3.651409945e-09 lua = -1.102674415e-14 wua = -1.169941157e-15 pua = 9.212818632e-21
+ ub = -8.051487260e-19 lub = 7.466843180e-24 wub = 8.536786732e-25 pub = -6.722378080e-30
+ uc = -6.821380085e-11 luc = 1.819443564e-16 wuc = 8.708731598e-18 puc = -6.857777784e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.321928268e-02 lu0 = -4.011701333e-08 wu0 = -4.586744968e-09 pu0 = 3.611878192e-14
+ a0 = 9.623533007e-01 la0 = -4.285908599e-07 wa0 = -1.908168637e-08 pa0 = 1.502606475e-13
+ keta = -7.160439798e-05 lketa = -6.386533375e-08 wketa = -6.775909406e-09 pketa = 5.335757621e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.626685010e-01 lags = -3.597756775e-07 wags = -4.176057083e-08 pags = 3.288477910e-13
+ b0 = 2.869435434e-07 lb0 = -2.259565627e-12 wb0 = -2.983627486e-13 pb0 = 2.349487300e-18
+ b1 = 9.463494026e-10 lb1 = -7.452123006e-15 wb1 = -9.840103234e-16 pb1 = 7.748687693e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.545664567e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 3.692110686e-07 wvoff = 3.806619356e-08 pvoff = -2.997560478e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '7.787032064e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.430654408e-05 wnfactor = -2.361338403e-06 pnfactor = 1.859459539e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 2.390451147e-02 ltvoff = -1.294608767e-07 wtvoff = -9.576639840e-09 ptvoff = 7.541220808e-14
+ cit = 1.567500000e-07 lcit = 3.813865645e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.716622884e-01 lpclm = 4.371927038e-06 wpclm = -2.587784236e-07 ppclm = 2.037776575e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 5.518791312e-03 lpdiblc2 = -1.638487482e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.260448608e+08 lpscbe1 = -1.045156920e+01 wpscbe1 = -1.723585164e+00 ppscbe1 = 1.357254373e-5
+ pscbe2 = 1.495053151e-08 lpscbe2 = 3.794886928e-16 wpscbe2 = 4.138093535e-17 ppscbe2 = -3.258583135e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.845482755e-04 lalpha0 = -9.473587494e-10 walpha0 = -6.038833331e-11 palpha0 = 4.755339695e-16
+ alpha1 = -4.028793582e-10 lalpha1 = 3.172513794e-15 walpha1 = 3.181925056e-16 palpha1 = -2.505638704e-21
+ beta0 = 1.800948224e+02 lbeta0 = -1.110754415e-03 wbeta0 = -1.103698784e-04 pbeta0 = 8.691186448e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.286240342e-07 lagidl = 2.343670220e-12 wagidl = 2.758983577e-13 pagidl = -2.172589208e-18
+ bgidl = 2.269601031e+09 lbgidl = -5.899658441e+03 wbgidl = -7.305699928e+02 pbgidl = 5.752946465e-3
+ cgidl = 4.446115856e+03 lcgidl = -2.398694392e-02 wcgidl = -2.252802939e-03 pcgidl = 1.773992203e-8
+ egidl = -1.732629844e+00 legidl = 2.561264870e-05 wegidl = 2.898483626e-06 pegidl = -2.282439916e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 1.474191273e-01 lkt1 = -7.592918686e-06 wkt1 = -8.592470420e-07 pkt1 = 6.766226757e-12
+ kt2 = -0.019032
+ at = 4.879756786e+05 lat = -2.652839965e+00 wat = -4.193459031e-01 pat = 3.302181248e-6
+ ute = -1.697232305e+00 lute = 1.111360449e-6
+ ua1 = 2.2096e-11
+ ub1 = -3.732379185e-18 lub1 = 5.163211310e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.67 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.564166162e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 2.273781170e-07 wvth0 = 1.324798710e-07 pvth0 = -1.940957865e-13
+ k1 = 7.249593021e-01 lk1 = -4.724807892e-08 wk1 = -1.133043617e-07 pk1 = 5.249056304e-15
+ k2 = -2.097029151e-02 lk2 = 2.032691772e-08 wk2 = 3.393877145e-08 pk2 = 3.631249432e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.040397055e+05 lvsat = 1.330520722e-01 wvsat = 3.298400555e-01 pvsat = -5.128089416e-7
+ ua = 1.137626284e-09 lua = -1.286837977e-15 wua = 1.169751432e-15 pua = 1.474457291e-22
+ ub = -5.367880817e-19 lub = 6.427053028e-24 wub = 6.586565747e-25 pub = -5.966745457e-30
+ uc = -1.441908912e-12 luc = -7.677001614e-17 wuc = -4.673064531e-17 puc = 1.462276319e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 9.993053255e-03 lu0 = 1.112933521e-08 wu0 = 8.550003932e-09 pu0 = -1.478086537e-14
+ a0 = 1.869742863e-01 la0 = 2.575692670e-06 wa0 = 6.463962910e-07 pa0 = -2.428200324e-12
+ keta = 3.056567038e-01 lketa = -1.248440237e-06 wketa = -2.256543593e-07 pketa = 9.014240180e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.250941926e+00 lags = 5.117399284e-06 wags = 8.582184185e-07 pags = -3.158210801e-12
+ b0 = -1.257537340e-07 lb0 = -6.605287557e-13 wb0 = 1.307582296e-13 pb0 = 6.868151580e-19
+ b1 = -8.551282568e-10 lb1 = -4.721176665e-16 wb1 = 8.891589409e-16 pb1 = 4.909060612e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-3.215452587e-03+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -2.172135321e-07 wvoff = -1.082257641e-07 pvoff = 2.670667715e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '-8.922628305e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 9.322251924e-06 wnfactor = 5.093381570e-06 pnfactor = -1.028946262e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -1.185842367e-02 ltvoff = 9.106191784e-09 wtvoff = 1.233034149e-08 ptvoff = -9.468581792e-15
+ cit = 2.190580279e-05 lcit = -4.613022348e-11 wcit = -9.403155419e-12 pcit = 3.643346598e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 3.326502231e-01 leta0 = -9.789184254e-07 weta0 = -1.847365935e-07 peta0 = 7.157804051e-13
+ etab = -1.330848348e-01 letab = 2.444285007e-07 wetab = -1.995155210e-09 petab = 7.730428375e-15
+ dsub = 1.006880630e+00 ldsub = -1.731483689e-06 wdsub = -1.722844542e-07 pdsub = 6.675333462e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.681793371e+00 lpclm = 1.293530093e-05 wpclm = 2.773729469e-06 ppclm = -9.711978505e-12
+ pdiblc1 = 8.502265248e-01 lpdiblc1 = -1.783193693e-06 wpdiblc1 = -4.794269295e-07 ppdiblc1 = 1.857587581e-12
+ pdiblc2 = 3.483154679e-03 lpdiblc2 = -8.497597119e-09 wpdiblc2 = -2.280433463e-09 ppdiblc2 = 8.835767494e-15
+ pdiblcb = -0.025
+ drout = -1.413331793e-01 ldrout = 2.717385537e-06 wdrout = 6.532244072e-07 pdrout = -2.530983288e-12
+ pscbe1 = 4.815713393e+07 lpscbe1 = 6.787922174e+02 wpscbe1 = 1.012526653e+02 ppscbe1 = -3.854192362e-4
+ pscbe2 = 1.455949168e-08 lpscbe2 = 1.894611616e-15 wpscbe2 = 6.991172876e-16 ppscbe2 = -2.874323584e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.362735909e-03 lalpha0 = 5.047748552e-09 walpha0 = 1.105321998e-09 palpha0 = -4.041127279e-15
+ alpha1 = 1.101869033e-09 lalpha1 = -2.657784321e-15 walpha1 = -9.442793336e-16 palpha1 = 2.385934684e-21
+ beta0 = -4.133476299e+02 lbeta0 = 1.188597711e-03 wbeta0 = 3.819025447e-04 pbeta0 = -1.038240086e-9
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.980422520e-07 lagidl = 1.077969027e-12 wagidl = 1.975961561e-14 pagidl = -1.180154038e-18
+ bgidl = -1.766712658e+09 lbgidl = 9.739442580e+03 wbgidl = 3.237998120e+03 pbgidl = -9.623667547e-3
+ cgidl = -1.709628086e+03 lcgidl = -1.358984407e-04 wcgidl = 1.950083002e-03 pcgidl = 1.455420157e-9
+ egidl = 6.463091431e+00 legidl = -6.142492957e-06 wegidl = -4.111565000e-06 pegidl = 4.336735245e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -2.642448653e+00 lkt1 = 3.216703014e-06 wkt1 = 1.608483443e-06 pkt1 = -2.795241779e-12
+ kt2 = -0.019032
+ at = -3.436518258e+05 lat = 5.693839638e-01 wat = 7.833816701e-01 pat = -1.357907007e-6
+ ute = -1.552796926e+00 lute = 5.517311276e-07 wute = 1.416313883e-07 pute = -5.487649772e-13
+ ua1 = -1.336349102e-09 lua1 = 5.263431393e-15 wua1 = 6.803232949e-16 pua1 = -2.635980639e-21
+ ub1 = -4.363120469e-18 lub1 = 7.607081489e-24 wub1 = 2.432365147e-24 pub1 = -9.424442001e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.68 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.924723990e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -7.995171263e-08 wvth0 = -9.776242920e-09 pvth0 = 7.257752460e-14
+ k1 = 6.896059835e-01 lk1 = 1.902525221e-08 wk1 = -1.024886547e-07 pk1 = -1.502606809e-14
+ k2 = -1.305601326e-02 lk2 = 5.490811722e-09 wk2 = 3.886884359e-08 pk2 = -5.610663812e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.685475856e+04 lvsat = 7.107170796e-03 wvsat = 3.763795723e-02 pvsat = 3.495311180e-8
+ ua = 3.055080055e-09 lua = -4.881296815e-15 wua = -8.079929975e-16 pua = 3.854925436e-21
+ ub = 7.599774430e-19 lub = 3.996136375e-24 wub = -8.576425227e-25 pub = -3.124291169e-30
+ uc = -7.911871300e-11 luc = 6.884292080e-17 wuc = 6.027858088e-17 puc = -5.437186348e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.255243979e-02 lu0 = -1.241449079e-08 wu0 = -4.292707187e-09 pu0 = 9.294080899e-15
+ a0 = 1.880524371e+00 la0 = -5.990363193e-07 wa0 = -9.013028515e-07 pa0 = 4.731164888e-13
+ keta = -4.475396235e-01 lketa = 1.635015986e-07 wketa = 3.209386003e-07 pketa = -1.232191441e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.576585638e+00 lags = -1.830838889e-07 wags = -9.036559676e-07 pags = 1.445989231e-13
+ b0 = -2.388331731e-07 lb0 = -4.485500392e-13 wb0 = 2.483377781e-13 pb0 = 4.664005365e-19
+ b1 = -1.282982596e-09 lb1 = 3.299380773e-16 wb1 = 1.334040171e-15 pb1 = -3.430682930e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.427791032e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 4.441248738e-08 wvoff = 5.295186116e-08 pvoff = -3.507680489e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.400437224e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.474043598e-06 wnfactor = -1.099382782e-06 pnfactor = 1.319493435e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -1.152340484e-02 ltvoff = 8.478165492e-09 wtvoff = 1.198199026e-08 ptvoff = -8.815562566e-15
+ cit = 4.376506056e-06 lcit = -1.326980383e-11 wcit = 4.441413023e-12 pcit = 1.048043798e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -3.993957024e-01 leta0 = 3.933748791e-07 weta0 = 3.793303798e-07 peta0 = -3.416195431e-13
+ etab = -1.418602834e-02 letab = 2.154079823e-08 wetab = 1.420243119e-08 petab = -2.263356710e-14
+ dsub = -9.106592846e-02 ldsub = 3.267269297e-07 wdsub = 3.214640620e-07 pdsub = -2.580476222e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.530545140e+00 lpclm = -4.334148843e-06 wpclm = -4.233137022e-06 ppclm = 3.423093419e-12
+ pdiblc1 = 1.378308749e-01 lpdiblc1 = -4.477368077e-07 wpdiblc1 = 3.228598737e-07 ppdiblc1 = 3.536207398e-13
+ pdiblc2 = -3.678778910e-03 lpdiblc2 = 4.928163587e-09 wpdiblc2 = 4.509287748e-09 ppdiblc2 = -3.892243888e-15
+ pdiblcb = -0.025
+ drout = -8.569112396e-03 ldrout = 2.468506017e-06 wdrout = 3.430957877e-07 pdrout = -1.949616178e-12
+ pscbe1 = 4.061302699e+08 lpscbe1 = 7.735776653e+00 wpscbe1 = -1.010889280e+02 ppscbe1 = -6.109685458e-6
+ pscbe2 = 1.684156675e-08 lpscbe2 = -2.383366308e-15 wpscbe2 = -1.838328973e-15 ppscbe2 = 1.882373177e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.223133010e-03 lalpha0 = -1.674321323e-09 walpha0 = -1.755821480e-09 palpha0 = 1.322372284e-15
+ alpha1 = -3.159184000e-10 walpha1 = 3.284906886e-16
+ beta0 = 2.403197680e+02 lbeta0 = -3.676719319e-05 wbeta0 = -1.874342035e-04 pbeta0 = 2.903858212e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.444895890e-06 lagidl = -1.259382803e-12 wagidl = -1.140185354e-12 pagidl = 9.942788034e-19
+ bgidl = 3.656480244e+09 lbgidl = -4.268748345e+02 wbgidl = -2.075568285e+03 pbgidl = 3.371440368e-4
+ cgidl = -1.904356087e+03 lcgidl = 2.291386691e-04 wcgidl = 3.289921468e-03 pcgidl = -1.056241030e-9
+ egidl = 8.122905745e+00 legidl = -9.253980869e-06 wegidl = -5.696981532e-06 pegidl = 7.308757074e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -8.420243340e-01 lkt1 = -1.583724135e-07 wkt1 = -1.560039006e-08 pkt1 = 2.492657740e-13
+ kt2 = -0.019032
+ at = -1.010637488e+05 lat = 1.146283547e-01 wat = 1.106202722e-01 pat = -9.674849005e-8
+ ute = -1.091146909e+00 lute = -3.136779934e-07 wute = -2.832627767e-07 pute = 2.477416245e-13
+ ua1 = 2.275182326e-09 lua1 = -1.506745422e-15 wua1 = -1.360646590e-15 pua1 = 1.190021507e-21
+ ub1 = 2.568576998e-18 lub1 = -5.387078582e-24 wub1 = -4.864730295e-24 pub1 = 4.254693116e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.69 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.508917816e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 5.860187939e-08 wvth0 = 9.832577431e-08 pvth0 = -2.196849967e-14
+ k1 = 9.822576657e-01 lk1 = -2.369279091e-07 wk1 = -3.336237827e-07 pk1 = 1.871247149e-13
+ k2 = -1.129682355e-01 lk2 = 9.287404125e-08 wk2 = 1.070336302e-07 pk2 = -6.522758619e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.906272476e+05 lvsat = 1.415965897e-01 wvsat = 2.192503523e-01 pvsat = -1.238850889e-7
+ ua = -8.642048819e-09 lua = 5.349012098e-15 wua = 8.428009998e-15 pua = -4.222882784e-21
+ ub = 1.028762302e-17 lub = -4.336742446e-24 wub = -7.947680351e-24 pub = 3.076655915e-30
+ uc = -5.062864152e-12 luc = 4.073675402e-18 wuc = 1.789567680e-18 puc = -3.217372538e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -2.353436102e-03 lu0 = 9.368188265e-09 wu0 = 1.603892151e-08 pu0 = -8.487961562e-15
+ a0 = 1.939538329e+00 la0 = -6.506499270e-07 wa0 = -9.479118395e-07 pa0 = 5.138807097e-13
+ keta = -5.806932352e-01 lketa = 2.799577473e-07 wketa = 4.328644693e-07 pketa = -2.211095090e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 2.652572021e-01 lags = 9.638039614e-07 wags = 1.320259860e-07 pags = -7.612085135e-13
+ b0 = -3.287167662e-06 lb0 = 2.217523305e-12 wb0 = 3.417983786e-12 pb0 = -2.305771862e-18
+ b1 = -3.960792505e-09 lb1 = 2.671950624e-15 wb1 = 4.118416203e-15 pb1 = -2.778283571e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-3.629792787e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -4.871594859e-08 wvoff = -3.114654522e-08 pvoff = 3.847566133e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.304897349e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.390484424e-06 wnfactor = -2.488118230e-06 pnfactor = 2.534081457e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -2.529027232e-02 ltvoff = 2.051866779e-08 wtvoff = 2.197441139e-08 ptvoff = -1.755493409e-14
+ cit = -8.094055816e-05 lcit = 6.134850053e-11 wcit = 7.182448907e-11 pcit = -4.845280033e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 5.093768088e-01 leta0 = -4.014375942e-07 weta0 = -3.737834427e-07 peta0 = 3.170538061e-13
+ etab = 5.685574834e-02 letab = -4.059233965e-08 wetab = -4.833271011e-08 petab = 3.205966749e-14
+ dsub = 8.816512678e-01 ldsub = -5.240115301e-07 wdsub = -4.467840888e-07 pdsub = 4.138622105e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.191983055e+00 lpclm = -1.414242443e-06 wpclm = -1.596354042e-06 ppclm = 1.116963025e-12
+ pdiblc1 = -2.182220839e+00 lpdiblc1 = 1.581380421e-06 wpdiblc1 = 2.155227437e-06 ppdiblc1 = -1.248967931e-12
+ pdiblc2 = -6.244912111e-02 lpdiblc2 = 5.632870488e-08 wpdiblc2 = 5.092586894e-08 ppdiblc2 = -4.448818580e-14
+ pdiblcb = -0.025
+ drout = 9.181619229e+00 ldrout = -5.569232706e-06 wdrout = -6.915278203e-06 pdrout = 4.398557715e-12
+ pscbe1 = -3.970616381e+08 lpscbe1 = 7.102074194e+02 wpscbe1 = 5.332688282e+02 ppscbe1 = -5.609189790e-4
+ pscbe2 = 2.722002529e-08 lpscbe2 = -1.146036615e-14 wpscbe2 = -1.003519402e-14 ppscbe2 = 9.051351343e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.948367573e-04 lalpha0 = -5.125934208e-10 walpha0 = -7.067384126e-10 palpha0 = 4.048442334e-16
+ alpha1 = -3.159184000e-10 walpha1 = 3.284906886e-16
+ beta0 = 2.334111594e+02 lbeta0 = -3.072492413e-05 wbeta0 = -1.819778120e-04 pbeta0 = 2.426642218e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.858310846e-07 lagidl = 3.417710093e-13 wagidl = 3.028218220e-13 pagidl = -2.677752732e-19
+ bgidl = -2.771044584e+08 lbgidl = 3.013438346e+03 wbgidl = 1.031161179e+03 pbgidl = -2.380001552e-3
+ cgidl = -3.744177492e+03 lcgidl = 1.838246470e-03 wcgidl = 3.742241018e-03 pcgidl = -1.451839709e-9
+ egidl = -3.329340165e+00 legidl = 7.621534033e-07 wegidl = 3.347956479e-06 pegidl = -6.019457093e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -9.059470176e-01 lkt1 = -1.024656345e-07 wkt1 = -5.688958436e-08 pkt1 = 2.853773034e-13
+ kt2 = -0.019032
+ at = -4.282927632e+04 lat = 6.369648507e-02 wat = 1.107999093e-01 pat = -9.690560066e-8
+ ute = -1.348610000e+00 lute = -8.850077400e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.70 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-9.299050203e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 4.444421021e-08 wvth0 = 1.633705933e-07 pvth0 = -6.584773458e-14
+ k1 = 2.150485169e-01 lk1 = 2.806313827e-07 wk1 = 2.519800171e-07 pk1 = -2.079236085e-13
+ k2 = 1.013767890e-01 lk2 = -5.172311222e-08 wk2 = -5.729514342e-08 pk2 = 4.562860450e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.282785567e+05 lvsat = 9.953616284e-02 wvsat = 1.609202742e-01 pvsat = -8.453561824e-8
+ ua = -7.089866449e-09 lua = 4.301909872e-15 wua = 9.220417866e-15 pua = -4.757441132e-21
+ ub = 1.867927265e-17 lub = -9.997749285e-24 wub = -1.881367411e-23 pub = 1.040685531e-29
+ uc = 9.143108392e-12 luc = -5.509673676e-18 wuc = -9.340104832e-18 puc = 4.290704538e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.660379578e-02 lu0 = -3.420360365e-09 wu0 = 1.157001823e-09 pu0 = 1.551381461e-15
+ a0 = 1.053076646e+00 la0 = -5.264287546e-08 wa0 = -3.807989218e-07 pa0 = 1.313063355e-13
+ keta = -5.992324220e-01 lketa = 2.924642828e-07 wketa = 5.234861416e-07 pketa = -2.822428892e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 5.736309113e+00 lags = -2.726967657e-06 wags = -5.166179022e-06 pags = 2.812960585e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-3.811344865e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.839107938e-07 wvoff = 3.003597289e-07 pvoff = -1.851584712e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '-1.878003614e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 2.455100566e-06 wnfactor = 5.525977452e-06 pnfactor = -2.872227490e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 9.152284876e-03 ltvoff = -2.716281294e-09 wtvoff = -5.194196601e-09 ptvoff = 7.730088631e-16
+ cit = -2.748371816e-05 lcit = 2.528651627e-11 wcit = 3.897542021e-11 pcit = -2.629281847e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -3.089567742e-01 leta0 = 1.506102409e-07 weta0 = 3.010732508e-07 peta0 = -1.382045193e-13
+ etab = -1.118725912e-02 letab = 5.309473177e-09 wetab = -2.727893766e-09 petab = 1.294658382e-15
+ dsub = -1.511509439e-01 ldsub = 1.727168419e-07 wdsub = 4.166073649e-07 pdsub = -1.685816642e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.980964394e+00 lpclm = -5.972892546e-07 wpclm = -7.309439242e-07 ppclm = 5.331573593e-13
+ pdiblc1 = 1.107147340e+00 lpdiblc1 = -6.376273524e-07 wpdiblc1 = -5.418643139e-07 ppdiblc1 = 5.704901641e-13
+ pdiblc2 = 2.762091489e-02 lpdiblc2 = -4.432541410e-09 wpdiblc2 = -2.492427538e-08 ppdiblc2 = 6.680321561e-15
+ pdiblcb = -0.025
+ drout = 4.274434259e+00 ldrout = -2.258845726e-06 wdrout = -4.114047273e-06 pdrout = 2.508847329e-12
+ pscbe1 = 1.869334997e+09 lpscbe1 = -8.187037504e+02 wpscbe1 = -1.485116929e+03 ppscbe1 = 8.006840528e-4
+ pscbe2 = -1.185982262e-09 lpscbe2 = 7.702326548e-15 wpscbe2 = 1.246370435e-14 ppscbe2 = -6.126405495e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.195229497e-04 lalpha0 = -1.919467262e-10 walpha0 = -3.955610143e-10 palpha0 = 1.949239605e-16
+ alpha1 = -1.065592763e-09 lalpha1 = 5.057303254e-16 walpha1 = 1.107999093e-15 palpha1 = -5.258563694e-22
+ beta0 = 5.292816288e+02 lbeta0 = -2.303191428e-04 wbeta0 = -5.028040822e-04 pbeta0 = 2.406958241e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.323281682e-06 lagidl = -8.111964630e-13 wagidl = -1.680740608e-12 pagidl = 1.070335942e-18
+ bgidl = 1.189584110e+10 lbgidl = -5.198430725e+03 wbgidl = -9.917777732e+03 pbgidl = 5.006152637e-3
+ cgidl = -6.974655772e+03 lcgidl = 4.017527118e-03 wcgidl = 6.657364360e-03 pcgidl = -3.418381915e-9
+ egidl = -1.224667412e+01 legidl = 6.777786891e-06 wegidl = 1.030913338e-05 pegidl = -5.297955648e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.588232997e+00 lkt1 = 3.578044870e-07 wkt1 = 7.344600123e-07 pkt1 = -2.484671346e-13
+ kt2 = -0.019032
+ at = 1.502892763e+05 lat = -6.658129054e-02 wat = -1.107999093e-01 pat = 5.258563694e-8
+ ute = -1.808697800e+00 lute = 2.218744559e-7
+ ua1 = 5.533492000e-10 lua1 = -6.403303200e-19
+ ub1 = -7.675544900e-18 lub1 = 2.755501450e-24
+ uc1 = 4.311053070e-10 luc1 = -3.644899601e-16 wuc1 = -5.618072970e-16 puc1 = 3.789952026e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.71 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-2.835309831e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.623249078e-07 wvth0 = -3.174839249e-07 pvth0 = 1.623658198e-13
+ k1 = 1.408911390e+00 lk1 = -2.859759371e-07 wk1 = -5.482666612e-07 pk1 = 1.718734650e-13
+ k2 = -8.518058405e-02 lk2 = 3.681701701e-08 wk2 = 1.717702635e-08 pk2 = 1.028411273e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.918101373e+05 lvsat = 1.771482510e-01 wvsat = 2.473402918e-01 pvsat = -1.255505586e-7
+ ua = 1.177553981e-08 lua = -4.651611939e-15 wua = -1.125318688e-14 pua = 4.959331681e-21
+ ub = -2.747177665e-17 lub = 1.190553871e-23 wub = 2.849282323e-23 pub = -1.204480833e-29
+ uc = 2.076809060e-11 luc = -1.102689023e-17 wuc = -1.201145892e-17 puc = 5.558529190e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -4.408388218e-03 lu0 = 6.552022162e-09 wu0 = 1.684822803e-08 pu0 = -5.895674497e-15
+ a0 = 1.318090465e+00 la0 = -1.784184342e-07 wa0 = -2.267071918e-08 pa0 = -3.866130950e-14
+ keta = -3.528588819e-01 lketa = 1.755354006e-07 wketa = 1.458976644e-07 pketa = -1.030393979e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 9.853252877e+00 lags = -4.680869168e-06 wags = -7.132389268e-06 pags = 3.746123968e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '6.188754533e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -2.906939236e-07 wvoff = -5.972801930e-07 pvoff = 2.408614357e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '1.525111438e+01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.674378834e-06 wnfactor = -8.500830321e-06 pnfactor = 3.784895480e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -6.329588158e-03 ltvoff = 4.631415647e-09 wtvoff = 6.581480448e-09 ptvoff = -4.815727464e-15
+ cit = 1.628689526e-04 lcit = -6.505486129e-11 wcit = -1.394771464e-10 pcit = 5.840076964e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.590369301e+00 leta0 = 7.587686262e-07 weta0 = 1.132578566e-06 peta0 = -5.328369420e-13
+ etab = 1.187988754e-01 letab = -5.638194625e-08 wetab = -8.089109553e-08 petab = 3.839091394e-14
+ dsub = -1.332732493e-01 ldsub = 1.642320880e-07 wdsub = 3.963622213e-07 pdsub = -1.589733190e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.743536160e+00 lpclm = -2.383005814e-06 wpclm = -3.040235682e-06 ppclm = 1.629147227e-12
+ pdiblc1 = -1.055603873e+00 lpdiblc1 = 3.888143733e-07 wpdiblc1 = 2.547108725e-06 ppdiblc1 = -8.955364403e-13
+ pdiblc2 = 9.823573802e-02 lpdiblc2 = -3.794633647e-08 wpdiblc2 = -7.151025796e-08 ppdiblc2 = 2.879002889e-14
+ pdiblcb = 3.091060653e+00 lpdiblcb = -1.478882386e-06 wpdiblcb = -2.461052239e-06 ppdiblcb = 1.168015393e-12
+ drout = -6.047992266e+00 ldrout = 2.640177903e-06 wdrout = 5.563204933e-06 pdrout = -2.083976568e-12
+ pscbe1 = -7.045694915e+09 lpscbe1 = 3.412369446e+03 wpscbe1 = 5.880580061e+03 ppscbe1 = -2.695075739e-3
+ pscbe2 = 1.572486853e-07 lpscbe2 = -6.749076669e-14 wpscbe2 = -1.135321084e-13 ppscbe2 = 5.367120725e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.392803618e-04 lalpha0 = -1.064035940e-10 walpha0 = -1.180394085e-10 palpha0 = 6.321220640e-17
+ alpha1 = 0.0
+ beta0 = 1.670725915e+02 lbeta0 = -5.841473370e-05 wbeta0 = -8.434327054e-05 pbeta0 = 4.209432282e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.049896290e-06 lagidl = -1.156047756e-12 wagidl = -1.729404383e-12 pagidl = 1.093431770e-18
+ bgidl = -6.293856091e+09 lbgidl = 3.434399560e+03 wbgidl = 6.216962215e+03 pbgidl = -2.651394942e-3
+ cgidl = 1.234027865e+04 lcgidl = -5.149340758e-03 wcgidl = -9.232808948e-03 pcgidl = 4.123094337e-9
+ egidl = 1.854575593e+01 legidl = -7.836300413e-06 wegidl = -1.382349612e-05 pegidl = 6.155390311e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -2.643624099e+00 lkt1 = 8.586931040e-07 wkt1 = 1.685531416e-06 pkt1 = -6.998456230e-13
+ kt2 = -0.019032
+ at = 9.105121306e+04 lat = -3.846690572e-02 wat = -4.922104479e-02 pat = 2.336030786e-8
+ ute = -3.553162726e+00 lute = 1.049797510e-06 wute = 1.831022866e-06 pute = -8.690034522e-13
+ ua1 = 5.52e-10
+ ub1 = -6.916664412e-18 lub1 = 2.395336770e-24 wub1 = 6.379047404e-24 pub1 = -3.027495898e-30
+ uc1 = -1.189810614e-09 luc1 = 4.047967360e-16 wuc1 = 1.123614594e-15 puc1 = -4.209060269e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.72 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.79342+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.57102
+ k2 = 0.0284341
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 180350.0
+ ua = 2.33476787e-9
+ ub = 6.10999999999999e-21
+ uc = -3.2639e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0188609
+ a0 = 0.87668
+ keta = -0.0076977
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1244
+ b0 = 9.3768e-8
+ b1 = 3.0925e-10
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.10903374+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.6003+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0030097
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.99495
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225600350.0
+ pscbe2 = 1.4994384e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.8978653e-5
+ alpha1 = 0.0
+ beta0 = 37.686511
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.15622e-7
+ bgidl = 1701900000.0
+ cgidl = 1200.0
+ egidl = 1.0890786
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.6891
+ kt2 = -0.019032
+ at = 351440.0
+ ute = -1.4104
+ ua1 = 2.2096e-11
+ ub1 = -2.3998e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.73 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.869956388e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.276816084e-7
+ k1 = 5.619445235e-01 lk1 = 1.803714652e-7
+ k2 = 3.148606463e-02 lk2 = -6.065657619e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.460989727e+05 lvsat = -1.306734533e+0
+ ua = 2.389660742e-09 lua = -1.090973873e-15
+ ub = -8.376543467e-20 lub = 1.786238314e-24 wub = 6.887662212e-41 pub = 1.401298464e-45
+ uc = -2.445625247e-11 luc = -1.626288342e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.934394109e-02 lu0 = -9.600248414e-9
+ a0 = 8.561756572e-01 la0 = 4.075156120e-7
+ keta = -7.379959890e-03 lketa = -6.314957590e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.292688783e-01 lags = -9.676700875e-8
+ b0 = 1.553001244e-07 lb0 = -1.222926360e-12
+ b1 = 5.121850042e-10 lb1 = -4.033252034e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.099220014e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.765384086e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.534658647e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 1.304595638e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 8.658285833e-05 ltvoff = 5.809578394e-8
+ cit = 1.328108333e-05 lcit = -6.521021882e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.593038174e+00 lpclm = -1.188676322e-5
+ pdiblc1 = 0.39
+ pdiblc2 = -1.195971040e-04 lpdiblc2 = 2.801517860e-08 ppdiblc2 = 2.524354897e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.261796187e+08 lpscbe1 = -1.151273371e+1
+ pscbe2 = 1.499153668e-08 lpscbe2 = 5.658942789e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.072433033e-05 lalpha0 = 5.903349124e-10
+ alpha1 = 0.0
+ beta0 = 3.679867151e+01 lbeta0 = 1.764545482e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.059446677e-08 lagidl = 6.961582120e-13
+ bgidl = 1.821003325e+09 lbgidl = -2.367130943e+3
+ cgidl = 1.068756667e+03 lcgidl = 2.608408753e-3
+ egidl = 8.063433181e-01 legidl = 5.619250633e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -6.052945695e-01 lkt1 = -1.665599409e-6
+ kt2 = -0.019032
+ at = 4.829130092e+05 lat = -2.612973468e+0
+ ute = -1.314789232e+00 lute = -1.900225776e-06 wute = 3.388131789e-21
+ ua1 = 2.2096e-11
+ ub1 = -1.955606938e-18 lub1 = -8.828159423e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.74 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.126930835e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 7.467548933e-8
+ k1 = 5.982464295e-01 lk1 = -1.054915237e-7
+ k2 = 1.927820612e-02 lk2 = 3.547542644e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.689691810e+04 lvsat = 7.642529089e-1
+ ua = 2.170089254e-09 lua = 6.380637651e-16
+ ub = 2.757363040e-19 lub = -1.044694077e-24
+ uc = -5.718724260e-11 luc = 9.511462079e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.741177674e-02 lu0 = 5.614773003e-9
+ a0 = 9.381930285e-01 la0 = -2.383383802e-7
+ keta = -8.650920330e-03 lketa = 3.693347491e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.097933651e-01 lags = 5.659486763e-8
+ b0 = -9.082837320e-08 lb0 = 7.152371076e-13
+ b1 = -2.995550125e-10 lb1 = 2.358875901e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.063689557e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.032497335e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.797224059e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -7.630019609e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 1.177905142e-02 ltvoff = -3.397772903e-08 wtvoff = -2.646977960e-23
+ cit = 1.567500000e-07 lcit = 3.813865645e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -7.993145222e-01 lpclm = 6.952057318e-06 wpclm = 4.235164736e-22 ppclm = -3.231174268e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 5.518791312e-03 lpdiblc2 = -1.638487482e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.238625439e+08 lpscbe1 = 6.733303519e+0
+ pscbe2 = 1.500292597e-08 lpscbe2 = -3.309672607e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.080876030e-04 lalpha0 = -3.452615376e-10
+ alpha1 = 0.0
+ beta0 = 4.035002948e+01 lbeta0 = -1.032006872e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.207045997e-07 lagidl = -4.071530408e-13
+ bgidl = 1.344590025e+09 lbgidl = 1.384433229e+3
+ cgidl = 1.593730000e+03 lcgidl = -1.525546258e-3
+ egidl = 1.937284446e+00 legidl = -3.286458369e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -9.405162915e-01 lkt1 = 9.741375630e-7
+ kt2 = -0.019032
+ at = -4.297902750e+04 lat = 1.528215964e+00 pat = -1.694065895e-21
+ ute = -1.697232305e+00 lute = 1.111360449e-6
+ ua1 = 2.2096e-11
+ ub1 = -3.732379185e-18 lub1 = 5.163211310e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.75 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.886772620e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.837621265e-8
+ k1 = 5.814990140e-01 lk1 = -4.060198764e-8
+ k2 = 2.200127513e-02 lk2 = 2.492462325e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.135871950e+05 lvsat = -5.162408357e-1
+ ua = 2.618706755e-09 lua = -1.100149605e-15
+ ub = 2.971697690e-19 lub = -1.127740181e-24 wub = 3.673419846e-40 pub = -1.751623080e-46
+ uc = -6.060990332e-11 luc = 1.083760620e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.081863851e-02 lu0 = -7.585453631e-9
+ a0 = 1.005408782e+00 la0 = -4.987725387e-7
+ keta = 1.994449549e-02 lketa = -1.071024506e-07 pketa = -5.048709793e-29
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.643088988e-01 lags = 1.118631499e-6
+ b0 = 3.980576440e-08 lb0 = 2.090820781e-13
+ b1 = 2.706801050e-10 lb1 = 1.494429152e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.402454757e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.209329911e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.556720920e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -3.705748497e-06 wnfactor = -1.355252716e-20
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 3.753635010e-03 ltvoff = -2.882450590e-9
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 9.874600000e-02 leta0 = -7.263325160e-08 weta0 = -2.117582368e-22
+ etab = -1.356110000e-01 letab = 2.542163806e-7
+ dsub = 7.887427130e-01 ldsub = -8.862865159e-07 wdsub = 1.694065895e-21
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.301634745e-01 lpclm = 6.384818719e-7
+ pdiblc1 = 2.432002427e-01 lpdiblc1 = 5.687903396e-7
+ pdiblc2 = 5.957844434e-04 lpdiblc2 = 2.689807596e-9
+ pdiblcb = -0.025
+ drout = 6.857467339e-01 ldrout = -4.872182953e-07 wdrout = -1.694065895e-21
+ pscbe1 = 1.763581697e+08 lpscbe1 = 1.907937516e+2
+ pscbe2 = 1.544467885e-08 lpscbe2 = -1.744712442e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.676725073e-05 lalpha0 = -6.892370075e-11
+ alpha1 = -9.373000000e-11 lalpha1 = 3.631662580e-16
+ beta0 = 7.019817776e+01 lbeta0 = -1.259697040e-4
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.230608842e-07 lagidl = -4.162827007e-13
+ bgidl = 2.333077820e+09 lbgidl = -2.445561581e+3
+ cgidl = 7.594690000e+02 lcgidl = 1.706881413e-3
+ egidl = 1.257234475e+00 legidl = -6.515367546e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -6.058677600e-01 lkt1 = -3.224916371e-7
+ kt2 = -0.019032
+ at = 6.482266720e+05 lat = -1.149929639e+0
+ ute = -1.373470380e+00 lute = -1.430875057e-7
+ ua1 = -4.749579392e-10 lua1 = 1.925885193e-15 wua1 = -1.972152263e-31
+ ub1 = -1.283381970e-18 lub1 = -4.325673299e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.76 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.048505864e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.194230127e-8
+ k1 = 0.55984
+ k2 = 3.615776294e-02 lk2 = -1.613128805e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.080053120e+04 lvsat = 5.136304421e-2
+ ua = 2.032039931e-09 lua = -3.839767925e-19
+ ub = -3.259264140e-19 lub = 4.031592368e-26
+ uc = -2.7970035e-12
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.711722970e-02 lu0 = -6.467926756e-10
+ a0 = 0.73934
+ keta = -4.118329820e-02 lketa = 7.487711406e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.43242187
+ b0 = 7.559964000e-08 lb0 = 1.419828789e-13
+ b1 = 4.061120200e-10 lb1 = -1.044377527e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.075734118+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.008454000e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -8.033673284e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 3.647589010e-03 ltvoff = -2.683656758e-9
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 8.089331940e-02 leta0 = -3.916661655e-8
+ etab = 3.796376220e-03 letab = -7.116686862e-9
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.1707598
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 278136550.0
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.250499886e-09 lagidl = -4.769542643e-16
+ bgidl = 1028500000.0
+ cgidl = 2.261177124e+03 lcgidl = -1.108220637e-3
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -8.617767638e-01 lkt1 = 1.572353814e-7
+ kt2 = -0.019032
+ at = 3.899808000e+04 lat = -7.869720768e-3
+ ute = -1.4498
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.77 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.263966280e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 3.078646925e-8
+ k1 = 0.55984
+ k2 = 2.255236760e-02 lk2 = 1.028614996e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.697652900e+04 lvsat = -1.526048346e-2
+ ua = 2.029073848e-09 lua = 2.210159329e-18
+ ub = 2.246696100e-19 lub = -4.412353589e-25
+ uc = -2.7970035e-12
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.795424020e-02 lu0 = -1.378842059e-9
+ a0 = 0.73934
+ keta = -0.032622
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.43242187
+ b0 = 1.040511620e-06 lb0 = -7.019291389e-13
+ b1 = 1.253739100e-09 lb1 = -8.457723969e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.075734118+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.154567100e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 8.180421543e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 2.532622950e-03 ltvoff = -1.708507442e-9
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.036111
+ etab = -0.0043407
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.1707598
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 278136550.0
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.413313420e-09 lagidl = 2.727416853e-15
+ bgidl = 1028500000.0
+ cgidl = 994.06
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -9.779777500e-01 lkt1 = 2.588647640e-7
+ kt2 = -0.019032
+ at = 9.746000000e+04 lat = -5.900051600e-2
+ ute = -1.348610000e+00 lute = -8.850077400e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.78 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.230533860e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -3.892888180e-8
+ k1 = 5.340929500e-01 lk1 = 1.736895993e-8
+ k2 = 2.883255802e-02 lk2 = 6.049533505e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.547060660e+04 lvsat = -7.498588212e-3
+ ua = 4.584563234e-09 lua = -1.721722980e-15
+ ub = -5.141655940e-18 lub = 3.178887857e-24 wub = -5.877471754e-39 pub = -1.401298464e-45
+ uc = -2.682862912e-12 luc = -7.699924073e-20
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.806873334e-02 lu0 = -1.456079131e-9
+ a0 = 5.709281900e-01 la0 = 1.136106070e-7
+ keta = 6.357942000e-02 lketa = -6.489747793e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -8.048471124e-01 lags = 8.346616555e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-8.340938640e-04+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.052755628e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.118711300e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.181569523e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 2.575654200e-03 ltvoff = -1.737536323e-9
+ cit = 2.186500000e-05 lcit = -8.004129000e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 7.224704400e-02 leta0 = -2.437737528e-8
+ etab = -1.464118110e-02 letab = 6.948704550e-9
+ dsub = 3.763363628e-01 ldsub = -4.073278837e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.055479935e+00 lpclm = 7.776779720e-8
+ pdiblc1 = 4.210659799e-01 lpdiblc1 = 8.469862052e-8
+ pdiblc2 = -3.936949901e-03 lpdiblc2 = 4.025745996e-9
+ pdiblcb = -0.025
+ drout = -9.345656259e-01 ldrout = 9.177306674e-7
+ pscbe1 = -1.104541685e+07 lpscbe1 = 1.950821548e+2
+ pscbe2 = 1.459493376e-08 lpscbe2 = -5.462017630e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -8.131652563e-05 lalpha0 = 5.485619565e-11 walpha0 = -5.219419293e-26 palpha0 = -3.541943154e-32
+ alpha1 = 3.373000000e-10 lalpha1 = -1.600825800e-16
+ beta0 = -1.073436291e+02 lbeta0 = 7.443781220e-05 wbeta0 = -2.710505431e-20 pbeta0 = -2.584939414e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.047876019e-07 lagidl = 5.440091119e-13 wagidl = -1.640830683e-28 pagidl = -3.731489267e-34
+ bgidl = -6.615506000e+08 lbgidl = 1.140108135e+3
+ cgidl = 1.454564380e+03 lcgidl = -3.106562547e-4
+ egidl = 8.062324272e-01 legidl = 6.978172551e-8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -6.582966430e-01 lkt1 = 4.320788917e-8
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.808697800e+00 lute = 2.218744559e-7
+ ua1 = 5.533492000e-10 lua1 = -6.403303200e-19
+ ub1 = -7.675544900e-18 lub1 = 2.755501450e-24
+ uc1 = -2.802268560e-10 luc1 = 1.153747171e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.79 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-6.855131720e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -5.674546737e-8
+ k1 = 7.147237000e-01 lk1 = -6.835839402e-8
+ k2 = -6.343189661e-02 lk2 = 4.983824367e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.135970880e+04 lvsat = 1.818244388e-2
+ ua = -2.472679832e-09 lua = 1.627644579e-15
+ ub = 8.604404080e-18 lub = -3.344992228e-24
+ uc = 5.559785013e-12 luc = -3.988959946e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.692399132e-02 lu0 = -9.127845685e-10
+ a0 = 1.289385940e+00 la0 = -2.273694411e-7
+ keta = -1.681305920e-01 lketa = 4.507209376e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 8.225800598e-01 lags = 6.228471960e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.373707077e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.427272065e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.487790280e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -8.821344069e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 2.003551600e-03 ltvoff = -1.466016429e-9
+ cit = -1.373000000e-05 lcit = 8.889258000e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.563552440e-01 leta0 = 8.411727060e-8
+ etab = 1.637863580e-02 letab = -7.773300551e-9
+ dsub = 3.685806741e-01 ldsub = -3.705193852e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.894142542e+00 lpclm = -3.202614761e-7
+ pdiblc1 = 2.169417177e+00 lpdiblc1 = -7.450688577e-7
+ pdiblc2 = 7.693043505e-03 lpdiblc2 = -1.493848874e-9
+ pdiblcb = -0.025
+ drout = 9.958582133e-01 ldrout = 1.551513313e-9
+ pscbe1 = 400000000.0
+ pscbe2 = 1.350003575e-08 lpscbe2 = 4.650184202e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.982479539e-05 lalpha0 = -2.636747531e-11
+ alpha1 = 0.0
+ beta0 = 6.028138144e+01 lbeta0 = -5.117017809e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.397886200e-07 lagidl = 2.284005951e-13
+ bgidl = 1.577749000e+09 lbgidl = 7.733654460e+1
+ cgidl = 6.501600000e+02 lcgidl = 7.111406400e-5
+ egidl = 1.043139921e+00 legidl = -4.265457116e-8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -5.094889340e-01 lkt1 = -2.741624952e-8
+ kt2 = -0.019032
+ at = 2.873000000e+04 lat = -8.889258000e-3
+ ute = -1.234813600e+00 lute = -5.049098544e-8
+ ua1 = 5.52e-10
+ ub1 = 1.160164800e-18 lub1 = -1.437926374e-24
+ uc1 = 2.328537120e-10 luc1 = -1.281333205e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.80 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.604296370e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = -2.440613859e-8
+ k1 = 5.188167327e-01 wk1 = 3.861976832e-8
+ k2 = 4.560035705e-02 wk2 = -1.269952830e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.326318546e+05 wvsat = -1.866371069e-1
+ ua = 3.565632057e-09 wua = -9.105884021e-16
+ ub = -1.414822211e-18 wub = 1.051199966e-24
+ uc = -1.774042234e-11 wuc = -1.102190816e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.953444859e-02 wu0 = -4.982885541e-10
+ a0 = 8.312423024e-01 wa0 = 3.361462691e-8
+ keta = -1.343529723e-02 wketa = 4.244651479e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.516368207e-01 wags = -2.014969101e-8
+ b0 = 2.089485401e-07 wb0 = -8.521010286e-14
+ b1 = -8.997671607e-10 wb1 = 8.944260594e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-8.744681044e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' wvoff = -1.596992414e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.543261839e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = 7.819926037e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 7.952014361e-03 wtvoff = -3.656304395e-9
+ cit = 2.627041256e-05 wcit = -1.203678613e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.491616770e+00 wpclm = -1.107228090e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.265862019e+08 wpscbe1 = -7.293292832e-1
+ pscbe2 = 1.498516181e-08 wpscbe2 = 6.822542275e-18
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.014387713e-05 walpha0 = -2.305590815e-11
+ alpha1 = -1.642128571e-10 walpha1 = 1.214840149e-16
+ beta0 = 9.464622176e+01 wbeta0 = -4.213856618e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.140183440e-07 wagidl = -7.279322171e-14
+ bgidl = 2.450053777e+09 wbgidl = -5.534811717e+2
+ cgidl = 8.715742857e+02 wcgidl = 2.429680297e-4
+ egidl = -4.067714573e-01 wegidl = 1.106623889e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 1.586488750e-01 wkt1 = -6.271612267e-7
+ kt2 = -0.019032
+ at = 8.516980480e+05 wat = -3.700889029e-1
+ ute = -1.353910777e+00 wute = -4.179050111e-8
+ ua1 = -1.101881891e-09 wua1 = 8.315143475e-16
+ ub1 = -1.176085789e-18 wub1 = -9.052988788e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.81 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.635527422e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 6.207046602e-08 wvth0 = -1.734296118e-08 pvth0 = -1.403778257e-13
+ k1 = 4.436740823e-01 lk1 = 1.493430120e-06 wk1 = 8.749599934e-08 pk1 = -9.713955409e-13
+ k2 = 6.930061527e-02 lk2 = -4.710331521e-07 wk2 = -2.797505331e-08 pk2 = 3.035949493e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.639323849e+05 lvsat = -4.597005521e+00 wvsat = -3.091114870e-01 pvsat = 2.434129316e-6
+ ua = 4.388214262e-09 lua = -1.634849228e-14 wua = -1.478521900e-15 pua = 1.128745109e-20
+ ub = -2.362790730e-18 lub = 1.884049513e-23 wub = 1.686013797e-24 pub = -1.261667098e-29
+ uc = 1.483395189e-11 luc = -6.474026581e-16 wuc = -2.906673602e-17 puc = 3.586337358e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.262902129e-02 lu0 = -6.150339463e-08 wu0 = -2.430289196e-09 pu0 = 3.839773996e-14
+ a0 = 7.508278238e-01 la0 = 1.598205596e-06 wa0 = 7.793590570e-08 pa0 = -8.808676873e-13
+ keta = -1.361852970e-02 lketa = 3.641672141e-09 wketa = 4.615268994e-09 pketa = -7.365874849e-15
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.766738165e-01 lags = -4.976002760e-07 wags = -3.506998363e-08 pags = 2.965348478e-13
+ b0 = 4.148704678e-07 lb0 = -4.092615944e-12 wb0 = -1.920291018e-13 pb0 = 2.122984875e-18
+ b1 = 7.867294732e-08 lb1 = -1.581475871e-12 wb1 = -5.782301932e-14 pb1 = 1.166985740e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-9.515752322e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.532473323e-07 wvoff = -1.092270193e-08 pvoff = -1.003115226e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.874352079e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 1.329431390e-05 wnfactor = 1.228288158e-06 pnfactor = -8.869945615e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 5.329868704e-03 ltvoff = 5.211409609e-08 wtvoff = -3.878961895e-09 ptvoff = 4.425228749e-15
+ cit = 3.753443144e-05 lcit = -2.238678697e-10 wcit = -1.794252992e-11 pcit = 1.173742955e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.071842353e+00 lpclm = -3.140635138e-05 wpclm = -1.833809417e-06 ppclm = 1.444051324e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 2.255652067e-03 lpdiblc2 = -1.919194857e-08 wpdiblc2 = -1.757199836e-09 ppdiblc2 = 3.492364386e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.281167043e+08 lpscbe1 = -3.041812267e+01 wpscbe1 = -1.433048157e+00 ppscbe1 = 1.398613113e-5
+ pscbe2 = 1.497763881e-08 lpscbe2 = 1.495165443e-16 wpscbe2 = 1.028158593e-17 ppscbe2 = -6.874710899e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.833522378e-05 lalpha0 = 1.559740739e-09 walpha0 = 1.302846853e-11 palpha0 = -7.171625527e-16
+ alpha1 = -1.642128571e-10 walpha1 = 1.214840149e-16
+ beta0 = 9.230043566e+01 lbeta0 = 4.662156035e-05 wbeta0 = -4.105998311e-05 pbeta0 = -2.143640696e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.299339791e-07 lagidl = -3.163168806e-13 wagidl = -1.104807738e-13 pagidl = 7.490250236e-19
+ bgidl = 2.822606773e+09 lbgidl = -7.404341769e+03 wbgidl = -7.409822243e+02 pbgidl = 3.726508420e-3
+ cgidl = 6.164078566e+02 lcgidl = 5.071330712e-03 wcgidl = 3.346458403e-04 pcgidl = -1.822059814e-9
+ egidl = -1.153794424e+00 legidl = 1.484678265e-05 wegidl = 1.450102061e-06 pegidl = -6.826491274e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 9.115312636e-01 lkt1 = -1.496323632e-05 wkt1 = -1.122141684e-06 pkt1 = 9.837538597e-12
+ kt2 = -0.019032
+ at = 1.311448726e+06 lat = -9.137360823e+00 wat = -6.129474091e-01 pat = 4.826715668e-6
+ ute = -1.221230839e+00 lute = -2.636960693e-06 wute = -6.921412445e-08 pute = 5.450335444e-13
+ ua1 = -1.839454915e-09 lua1 = 1.465896884e-14 wua1 = 1.377167921e-15 pua1 = -1.084464651e-20
+ ub1 = 7.112893387e-20 lub1 = -2.478789372e-23 wub1 = -1.499371091e-24 pub1 = 1.180694760e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.82 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-8.071624708e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 4.054796353e-07 wvth0 = -4.091525131e-09 pvth0 = -2.447275840e-13
+ k1 = 7.246160897e-01 lk1 = -7.188758111e-07 wk1 = -9.348776913e-08 pk1 = 4.537792423e-13
+ k2 = -2.424242196e-02 lk2 = 2.655808489e-07 wk2 = 3.219638657e-08 pk2 = -1.702310711e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.125266663e+05 lvsat = 1.517298924e+00 wvsat = 7.074650519e-02 pvsat = -5.571004297e-7
+ ua = 1.940719278e-09 lua = 2.924551710e-15 wua = 1.696869905e-16 pua = -1.691534636e-21
+ ub = 7.943823297e-19 lub = -6.020979844e-24 wub = -3.836922552e-25 pub = 3.681436305e-30
+ uc = -9.278856738e-11 luc = 2.000816322e-16 wuc = 2.633771767e-17 puc = -7.765417516e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.397352723e-02 lu0 = 6.655158931e-09 wu0 = 2.543603231e-09 pu0 = -7.696733482e-16
+ a0 = 9.224081144e-01 la0 = 2.470794400e-07 wa0 = 1.167761631e-08 pa0 = -3.591101617e-13
+ keta = -1.424735342e-02 lketa = 8.593407389e-09 wketa = 4.140218815e-09 pketa = -3.625044713e-15
+ a1 = 0.0
+ a2 = 0.5
+ ags = 8.770045262e-02 lags = 2.030293749e-07 wags = 1.634424827e-08 pags = -1.083316628e-13
+ b0 = -3.404782397e-07 lb0 = 1.855452988e-12 wb0 = 1.846899726e-13 pb0 = -8.435271477e-19
+ b1 = -2.303445928e-07 lb1 = 8.519136499e-13 wb1 = 1.701863988e-13 pb1 = -6.284972236e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.094621570e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 2.658906015e-07 wvoff = 2.288337973e-09 pvoff = -2.043431774e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.847720095e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.245169874e-06 wnfactor = -3.735676523e-08 pnfactor = 1.096501894e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 1.951416253e-02 ltvoff = -5.958154406e-08 wtvoff = -5.722404253e-09 ptvoff = 1.894159994e-14
+ cit = 2.854518268e-07 lcit = 6.945294517e-11 wcit = -9.521309665e-14 pcit = -2.316618554e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -3.202563950e-01 lpclm = 3.179669422e-06 wpclm = -3.544052862e-07 ppclm = 2.790797475e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -1.606956202e-03 lpdiblc2 = 1.122454650e-08 wpdiblc2 = 5.271599508e-09 ppdiblc2 = -2.042533945e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.219969853e+08 lpscbe1 = 1.777221658e+01 wpscbe1 = 1.380132812e+00 ppscbe1 = -8.166543725e-6
+ pscbe2 = 1.500774829e-08 lpscbe2 = -8.758358843e-17 wpscbe2 = -3.567532989e-18 ppscbe2 = 4.030916283e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.206713007e-04 lalpha0 = -1.188546039e-09 walpha0 = -1.572685692e-10 palpha0 = 6.238585007e-16
+ alpha1 = -3.232776412e-10 lalpha1 = 1.252571549e-15 walpha1 = 2.391595059e-16 palpha1 = -9.266474214e-22
+ beta0 = 1.557077293e+02 lbeta0 = -4.526855143e-04 wbeta0 = -8.534116491e-05 pbeta0 = 3.272601872e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.107913390e-07 lagidl = -9.530362474e-13 wagidl = -6.664580941e-14 pagidl = 4.038422127e-19
+ bgidl = 1.872799261e+09 lbgidl = 7.501246818e+01 wbgidl = -3.907670796e+02 pbgidl = 9.687042413e-4
+ cgidl = 1.318944005e+03 lcgidl = -4.608604416e-04 wcgidl = 2.032855800e-04 pcgidl = -7.876503082e-10
+ egidl = 7.672350385e-01 legidl = -2.805559554e-07 wegidl = 8.655978711e-07 pegidl = -2.223754582e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.192929769e+00 lkt1 = 1.608552527e-06 wkt1 = 1.867344810e-07 pkt1 = -4.693376525e-13
+ kt2 = -0.019032
+ at = -2.526105064e+05 lat = 3.178980008e+00 wat = 1.550845296e-01 pat = -1.221228637e-6
+ ute = -1.748133036e+00 lute = 1.512183345e-06 wute = 3.765615712e-08 pute = -2.965271748e-13
+ ua1 = 2.2096e-11
+ ub1 = -3.732379185e-18 lub1 = 5.163211310e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.83 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-7.477103795e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.751265623e-07 wvth0 = -3.030713580e-08 pvth0 = -1.431525789e-13
+ k1 = 5.681835353e-01 lk1 = -1.127622359e-07 wk1 = 9.850737868e-09 pk1 = 5.338386305e-14
+ k2 = 2.612820761e-02 lk2 = 7.041480756e-08 wk2 = -3.053088145e-09 pk2 = -3.365345639e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.474505241e+05 lvsat = -1.427308698e+00 wvsat = -2.469907554e-01 pvsat = 6.740043602e-7
+ ua = 3.205428287e-09 lua = -1.975689816e-15 wua = -4.340542426e-16 pua = 6.477211461e-22
+ ub = 4.947551235e-19 lub = -4.860044270e-24 wub = -1.461728549e-25 pub = 2.761143636e-30
+ uc = -9.048780653e-11 luc = 1.911671042e-16 wuc = 2.210355329e-17 puc = -6.124848185e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.141499907e-02 lu0 = -2.217756784e-08 wu0 = -4.411851533e-10 pu0 = 1.079518772e-14
+ a0 = 1.434036824e+00 la0 = -1.735277157e-06 wa0 = -3.170973108e-07 pa0 = 9.147611707e-13
+ keta = 5.494013728e-02 lketa = -2.594804441e-07 wketa = -2.588963581e-08 pketa = 1.127286300e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -6.455450534e-01 lags = 3.044062412e-06 wags = 3.560165822e-07 pags = -1.424426088e-12
+ b0 = -2.713646221e-09 lb0 = 5.467502945e-13 wb0 = 3.145568990e-14 pb0 = -2.498055959e-19
+ b1 = 7.758929642e-08 lb1 = -3.412069971e-13 wb1 = -5.720000308e-14 pb1 = 2.525341289e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.201780836e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 3.074105306e-07 wvoff = -1.484577642e-08 pvoff = -1.379553377e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.851434499e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.259561702e-06 wnfactor = 5.217680733e-07 pnfactor = -1.069883206e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 2.526163920e-03 ltvoff = 6.240155346e-09 wtvoff = 9.080782022e-10 ptvoff = -6.748867381e-15
+ cit = 1.821064286e-05 wcit = -6.074200743e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 7.605878573e-01 leta0 = -2.637005712e-06 weta0 = -4.896279587e-07 peta0 = 1.897112489e-12
+ etab = -1.761741052e+00 letab = 6.554819879e-06 wetab = 1.203004508e-06 petab = -4.661161266e-12
+ dsub = 7.026175246e-01 ldsub = -5.525858607e-07 wdsub = 6.371506991e-08 pdsub = -2.468704099e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 9.526035596e-01 lpclm = -1.752153758e-06 wpclm = -9.058068523e-08 ppclm = 1.768582676e-12
+ pdiblc1 = 2.998208906e-01 lpdiblc1 = 3.494079774e-07 wpdiblc1 = -4.188772880e-08 ppdiblc1 = 1.622981940e-13
+ pdiblc2 = -5.442067568e-04 lpdiblc2 = 7.106817500e-09 wpdiblc2 = 8.433609299e-10 ppdiblc2 = -3.267686259e-15
+ pdiblcb = -0.025
+ drout = 5.078815216e-01 ldrout = 2.019382564e-07 wdrout = 1.315839726e-07 pdrout = -5.098352603e-13
+ pscbe1 = 2.008949618e+08 lpscbe1 = 9.953411689e+01 wpscbe1 = -1.815222059e+01 ppscbe1 = 6.751351275e-5
+ pscbe2 = 1.577727376e-08 lpscbe2 = -3.069186963e-15 wpscbe2 = -2.460523805e-16 ppscbe2 = 9.798409528e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.584328931e-05 lalpha0 = -8.495142581e-11 walpha0 = 6.835429613e-13 palpha0 = 1.185724689e-17
+ alpha1 = -2.476467110e-10 lalpha1 = 9.595319464e-16 walpha1 = 1.138669671e-16 palpha1 = -4.411889508e-22
+ beta0 = 1.221679331e+02 lbeta0 = -3.227322198e-04 wbeta0 = -3.844701710e-05 pbeta0 = 1.455641221e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.335766006e-07 lagidl = -1.428780022e-12 wagidl = -1.557386849e-13 pagidl = 7.490414681e-19
+ bgidl = 3.533512365e+09 lbgidl = -6.359586526e+03 wbgidl = -8.880766745e+02 pbgidl = 2.895579998e-3
+ cgidl = -3.781956298e+01 lcgidl = 4.796055679e-03 wcgidl = 5.898308897e-04 pcgidl = -2.285358765e-9
+ egidl = 1.365261907e+00 legidl = -2.597670861e-06 wegidl = -7.991826195e-08 pegidl = 1.439742227e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -8.302542482e-01 lkt1 = 2.033299541e-07 wkt1 = 1.660002265e-07 pkt1 = -3.890007099e-13
+ kt2 = -0.019032
+ at = 1.297133363e+06 lat = -2.825657587e+00 wat = -4.800585741e-01 pat = 1.239696833e-6
+ ute = -1.118060041e+00 lute = -9.290974830e-07 wute = -1.889515474e-07 pute = 5.814870372e-13
+ ua1 = -4.749579392e-10 lua1 = 1.925885193e-15 wua1 = 6.162975822e-33 pua1 = 1.175494351e-38
+ ub1 = -6.872625483e-19 lub1 = -6.635397610e-24 wub1 = -4.410067637e-25 pub1 = 1.708724807e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.84 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-6.085333631e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -8.577467274e-08 wvth0 = -1.452346966e-07 pvth0 = 7.229062650e-14
+ k1 = 4.950829183e-01 lk1 = 2.427218080e-08 wk1 = 4.790703005e-08 pk1 = -1.795646227e-14
+ k2 = 7.633295128e-02 lk2 = -2.369900491e-08 wk2 = -2.972144363e-08 pk2 = 1.633904280e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.456284455e+05 lvsat = 2.468571384e-01 wvsat = 1.897051312e-01 pvsat = -1.446257489e-7
+ ua = 1.870805342e-09 lua = 5.261943568e-16 wua = 1.192807041e-16 pua = -3.895605449e-22
+ ub = -2.148790005e-18 lub = 9.554542839e-26 wub = 1.348547193e-24 pub = -4.085856666e-32
+ uc = 2.183214270e-11 luc = -1.938787264e-17 wuc = -1.822054384e-17 puc = 1.434307063e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 8.116056594e-03 lu0 = 2.752629715e-09 wu0 = 6.659031859e-09 pu0 = -2.514879087e-15
+ a0 = 1.541575819e-01 la0 = 6.639844695e-07 wa0 = 4.329156122e-07 pa0 = -4.912130546e-13
+ keta = -9.919594011e-02 lketa = 2.946304660e-08 wketa = 4.291752043e-08 pketa = -1.625726508e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.018694604e+00 lags = -7.572124994e-08 wags = -4.337222238e-07 pags = 5.601827782e-14
+ b0 = 7.993566900e-08 lb0 = 3.918158882e-13 wb0 = -3.207776909e-15 pb0 = -1.848254610e-19
+ b1 = -1.946639869e-07 lb1 = 1.691590078e-13 wb1 = 1.443120789e-13 pb1 = -1.252204200e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '8.319962512e-02+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -7.384132217e-08 wvoff = -1.175785474e-07 pvoff = 5.462751477e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.303850203e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.233060181e-06 wnfactor = -2.185329294e-07 pnfactor = 3.178850539e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 9.377589538e-03 ltvoff = -6.603527117e-09 wtvoff = -4.239031471e-09 ptvoff = 2.899904412e-15
+ cit = 1.821064286e-05 wcit = -6.074200743e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -8.818302658e-01 leta0 = 4.418713016e-07 weta0 = 7.122190574e-07 peta0 = -3.558699277e-13
+ etab = 3.261181120e+00 letab = -2.861150024e-06 wetab = -2.409800204e-06 petab = 2.111402447e-12
+ dsub = 4.197837131e-01 ldsub = -2.238559764e-08 wdsub = -7.681154135e-08 pdsub = 1.656077559e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.274633399e+00 lpclm = 2.423024644e-06 wpclm = 1.809092107e-06 ppclm = -1.792543940e-12
+ pdiblc1 = 2.523648661e-01 lpdiblc1 = 4.383690409e-07 wpdiblc1 = 2.176886379e-07 ppdiblc1 = -3.243036630e-13
+ pdiblc2 = 3.078269865e-03 lpdiblc2 = 3.161228242e-10 wpdiblc2 = -7.750215827e-10 ppdiblc2 = -2.338664009e-16
+ pdiblcb = -0.025
+ drout = 1.427978215e+00 ldrout = -1.522875006e-06 wdrout = -7.413767112e-07 pdrout = 1.126616838e-12
+ pscbe1 = 2.771708354e+08 lpscbe1 = -4.345263591e+01 wpscbe1 = 7.144317738e-01 ppscbe1 = 3.214608624e-5
+ pscbe2 = 1.434404927e-08 lpscbe2 = -3.824643315e-16 wpscbe2 = 1.257044585e-16 ppscbe2 = 2.829455826e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.630807725e-06 lalpha0 = -1.282788351e-11 walpha0 = 1.946335011e-12 palpha0 = 9.490016909e-18
+ alpha1 = 2.642128571e-10 walpha1 = -1.214840149e-16
+ beta0 = -4.289798735e+01 lbeta0 = -1.329964534e-05 wbeta0 = 3.395514745e-05 pbeta0 = 9.839024423e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -4.161300340e-07 lagidl = 1.640800353e-13 wagidl = 3.087764494e-13 pagidl = -1.217386027e-19
+ bgidl = 4.511179773e+08 lbgidl = -5.813300069e+02 wbgidl = 4.271449109e+02 pbgidl = 4.300656138e-4
+ cgidl = 3.864285312e+03 lcgidl = -2.518830119e-03 wcgidl = -1.185973025e-03 pcgidl = 1.043563253e-9
+ egidl = -1.043567258e+00 legidl = 1.917920292e-06 wegidl = 1.445000114e-06 pegidl = -1.418869760e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -6.866934015e-01 lkt1 = -6.578920929e-08 wkt1 = -1.295259711e-07 pkt1 = 1.649927001e-13
+ kt2 = -0.019032
+ at = -4.490134986e+05 lat = 4.476693188e-01 wat = 3.610290138e-01 pat = -3.370059593e-7
+ ute = -1.757017755e+00 lute = 2.686926487e-07 wute = 2.272784664e-07 pute = -1.987777467e-13
+ ua1 = 5.524e-10
+ ub1 = -3.784975918e-18 lub1 = -8.284241282e-25 wub1 = 1.435765876e-25 pub1 = 6.128648563e-31
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.85 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.018191635e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 2.725124519e-07 wvth0 = 1.418891790e-07 pvth0 = -1.788279150e-13
+ k1 = 2.087157100e-01 lk1 = 2.747289412e-07 wk1 = 2.597603453e-07 pk1 = -2.032433718e-13
+ k2 = 1.496279473e-01 lk2 = -8.780280843e-08 wk2 = -9.401000556e-08 pk2 = 7.256581906e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.544260090e+04 lvsat = 6.302859876e-02 wvsat = 9.056518263e-02 pvsat = -5.791794988e-8
+ ua = 1.378690597e-09 lua = 9.565979128e-16 wua = 4.811509277e-16 pua = -7.060522425e-22
+ ub = -2.084927034e-18 lub = 3.969087389e-26 wub = 1.708630359e-24 pub = -3.557873033e-31
+ uc = -6.648391153e-13 luc = 2.879876558e-19 wuc = -1.577366683e-18 puc = -2.130521158e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.394964857e-03 lu0 = 6.007096548e-09 wu0 = 1.003109766e-08 pu0 = -5.464087837e-15
+ a0 = 1.643952427e+00 la0 = -6.389901023e-07 wa0 = -6.692286553e-07 pa0 = 4.727223217e-13
+ keta = -1.598406619e-01 lketa = 8.250292026e-08 wketa = 9.411585718e-08 pketa = -6.103533040e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 2.470985405e+00 lags = -1.345894784e-06 wags = -1.508121149e-06 pags = 9.956875779e-13
+ b0 = 2.308638122e-06 lb0 = -1.557407277e-12 wb0 = -9.381549133e-13 pb0 = 6.328793045e-19
+ b1 = -5.470575747e-09 lb1 = 3.690450399e-15 wb1 = 4.974621226e-15 pb1 = -3.355879479e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-1.153651976e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.007909088e-06 wvoff = 7.974393198e-07 pvoff = -7.456471119e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '1.511379504e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 1.209234692e-06 wnfactor = 4.758276107e-07 pnfactor = -2.894026745e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = -1.238095564e-02 ltvoff = 1.242649649e-08 wtvoff = 1.103300578e-08 ptvoff = -1.045701937e-14
+ cit = 1.821064286e-05 wcit = -6.074200743e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 7.453559857e-01 leta0 = -9.812657940e-07 weta0 = -5.246966035e-07 peta0 = 7.259365093e-13
+ etab = -5.955817675e-03 letab = -3.712058353e-09 wetab = 1.194857595e-09 petab = 2.746165921e-15
+ dsub = 1.506860750e+00 ldsub = -9.731431745e-07 wdsub = -8.810267853e-07 pdsub = 7.199274279e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.617412977e+00 lpclm = -1.063591165e-07 wpclm = -3.304322341e-07 ppclm = 7.868404895e-14
+ pdiblc1 = 6.487935858e-01 lpdiblc1 = 9.165248261e-08 wpdiblc1 = -7.558774327e-08 ppdiblc1 = -6.780414002e-14
+ pdiblc2 = 3.290184241e-02 lpdiblc2 = -2.576757373e-08 wpdiblc2 = -2.283838126e-08 ppdiblc2 = 1.906274797e-14
+ pdiblcb = -0.025
+ drout = -2.335481063e+00 ldrout = 1.768646479e-06 wdrout = 2.042815409e-06 pdrout = -1.308437590e-12
+ pscbe1 = 2.271135937e+08 lpscbe1 = 3.274277005e-01 wpscbe1 = 3.774657897e+01 ppscbe1 = -2.422297031e-7
+ pscbe2 = 1.145298702e-08 lpscbe2 = 2.146058714e-15 wpscbe2 = 2.264500748e-15 ppscbe2 = -1.587645652e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -7.564427703e-05 lalpha0 = 5.102969674e-11 walpha0 = 5.596140755e-11 palpha0 = -3.775156553e-17
+ alpha1 = 8.181028243e-10 lalpha1 = -4.844321653e-16 walpha1 = -5.312495970e-16 palpha1 = 3.583809781e-22
+ beta0 = -2.642101254e+02 lbeta0 = 1.802599506e-04 wbeta0 = 1.976809819e-04 pbeta0 = -1.333555904e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.857215868e-06 lagidl = -2.698788290e-12 wagidl = -2.115542230e-12 pagidl = 1.998570514e-18
+ bgidl = -1.266898348e+09 lbgidl = 9.212470708e+02 wbgidl = 1.698126516e+03 pbgidl = -6.815348980e-4
+ cgidl = 2.728410918e+04 lcgidl = -2.300180807e-02 wcgidl = -1.944927322e-02 pcgidl = 1.701664560e-8
+ egidl = 7.996957227e+00 legidl = -5.988922422e-06 wegidl = -5.243143738e-06 pegidl = 4.430580852e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -6.891749787e-01 lkt1 = -6.361882187e-08 wkt1 = -2.136551350e-07 pkt1 = 2.385720669e-13
+ kt2 = -0.019032
+ at = 2.410805649e+05 lat = -1.558869491e-01 wat = -1.062499194e-01 pat = 7.167619563e-8
+ ute = -1.348610000e+00 lute = -8.850077400e-8
+ ua1 = 5.524e-10
+ ub1 = -4.732179357e-18 wub1 = 8.443139033e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.86 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.841331924e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.901433735e-07 wvth0 = -3.986910035e-07 pvth0 = 1.858474761e-13
+ k1 = 5.822784973e-01 lk1 = 2.272348481e-08 wk1 = -3.564747518e-08 pk1 = -3.961256087e-15
+ k2 = 1.146295632e-02 lk2 = 5.403294480e-09 wk2 = 1.284996185e-08 pk2 = 4.780850453e-16
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.072378449e+05 lvsat = -3.322363000e-02 wvsat = -2.350127585e-02 pvsat = 1.903128302e-8
+ ua = 8.006101065e-09 lua = -3.514253189e-15 wua = -2.531240001e-15 pua = 1.326106678e-21
+ ub = -1.215456639e-17 lub = 6.832669580e-24 wub = 5.188123096e-24 pub = -2.703053103e-30
+ uc = -1.126486252e-12 luc = 5.994148145e-19 wuc = -1.151401227e-18 puc = -5.004084124e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.495383126e-02 lu0 = -1.115914728e-09 wu0 = 2.304392099e-09 pu0 = -2.516522651e-16
+ a0 = -2.619971856e-01 la0 = 6.467635066e-07 wa0 = 6.161948611e-07 pa0 = -3.944243825e-13
+ keta = 2.578804530e-01 lketa = -1.992917438e-07 wketa = -1.437431270e-07 pketa = 9.942434033e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = -2.690000976e+00 lags = 2.135706629e-06 wags = 1.394629288e-06 pags = -9.625078670e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '1.387059142e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -7.060546322e-07 wvoff = -1.026757865e-06 pvoff = 4.849563087e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.256629411e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.317310895e-06 wnfactor = -1.020312667e-07 pnfactor = 1.004209242e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 2.495981661e-02 ltvoff = -1.276358846e-08 wtvoff = -1.655971381e-08 ptvoff = 8.157029269e-15
+ cit = 6.904335386e-05 lcit = -3.429174684e-11 wcit = -3.490235747e-11 pcit = 1.944747453e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -2.155105805e+00 leta0 = 9.753857303e-07 weta0 = 1.647786729e-06 peta0 = -7.396207465e-13
+ etab = -1.785280447e-01 letab = 1.127051660e-07 wetab = 1.212428461e-07 petab = -7.823820713e-14
+ dsub = -4.580615905e-01 ldsub = 3.523934366e-07 wdsub = 6.172842682e-07 pdsub = -2.908332088e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.564235730e+00 lpclm = -7.048574508e-08 wpclm = -3.763755021e-07 ppclm = 1.096773776e-13
+ pdiblc1 = 2.676812648e-01 lpdiblc1 = 3.487508544e-07 wpdiblc1 = 1.134733987e-07 ppdiblc1 = -1.953447864e-13
+ pdiblc2 = -3.373360724e-02 lpdiblc2 = 1.918470061e-08 wpdiblc2 = 2.204344791e-08 ppdiblc2 = -1.121453399e-14
+ pdiblcb = -0.025
+ drout = -2.500905813e+00 ldrout = 1.880242016e-06 wdrout = 1.158772205e-06 pdrout = -7.120620454e-13
+ pscbe1 = -2.399248548e+08 lpscbe1 = 3.153915650e+02 wpscbe1 = 1.693240927e+02 ppscbe1 = -8.900442043e-5
+ pscbe2 = 1.236987844e-08 lpscbe2 = 1.527523762e-15 wpscbe2 = 1.646087029e-15 ppscbe2 = -1.170463757e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.375038343e-04 lalpha0 = 9.276015409e-11 walpha0 = 4.156714622e-11 palpha0 = -2.804119684e-17
+ alpha1 = 3.373000000e-10 lalpha1 = -1.600825800e-16
+ beta0 = -1.245301003e+02 lbeta0 = 8.603180569e-05 wbeta0 = 1.271448267e-05 pbeta0 = -8.577190011e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.883518583e-06 lagidl = 1.173911170e-12 wagidl = 1.537836865e-12 pagidl = -4.659990233e-19
+ bgidl = -4.419883131e+09 lbgidl = 3.048250605e+03 wbgidl = 2.780399373e+03 pbgidl = -1.411636167e-3
+ cgidl = -2.055973837e+04 lcgidl = 9.273651484e-03 wcgidl = 1.628609312e-02 pcgidl = -7.090432528e-9
+ egidl = -3.729696459e+00 legidl = 1.921878154e-06 wegidl = 3.355662046e-06 pegidl = -1.370173529e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.349333415e+00 lkt1 = 3.817240591e-07 wkt1 = 5.112262396e-07 pkt1 = -2.504329085e-13
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.419020690e+00 lute = -4.100172253e-08 wute = -2.882815673e-07 pute = 1.944747453e-13
+ ua1 = 5.533492000e-10 lua1 = -6.403303200e-19
+ ub1 = -1.152508017e-17 lub1 = 4.582490889e-24 wub1 = 2.847870796e-24 pub1 = -1.351599480e-30
+ uc1 = -5.610749427e-10 luc1 = 3.048348364e-16 wuc1 = 2.077702912e-16 puc1 = -1.401618384e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.87 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 6.27e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.9898e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.1045e-08+MC_MM_SWITCH*GAU*(1.1045e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-4.260212896e-01+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.753432825e-07 wvth0 = -1.919710566e-07 pvth0 = 8.773818927e-14
+ k1 = 8.257022010e-01 lk1 = -9.280540497e-08 wk1 = -8.210145115e-08 pk1 = 1.808580091e-14
+ k2 = -9.392889550e-02 lk2 = 5.542226735e-08 wk2 = 2.256155779e-08 pk2 = -4.131038386e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.562912187e+04 lvsat = 3.458103245e-02 wvsat = 4.216010898e-02 pvsat = -1.213161023e-8
+ ua = -2.015020126e-10 lua = 3.810752320e-16 wua = -1.680208266e-15 pua = 9.222070166e-22
+ ub = 2.579848447e-18 lub = -1.602836994e-25 wub = 4.456942159e-24 pub = -2.356034631e-30
+ uc = 7.667866730e-12 luc = -3.574385111e-18 wuc = -1.559550422e-18 puc = -3.067008045e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.369354828e-02 lu0 = -5.177844271e-10 wu0 = 2.389868836e-09 pu0 = -2.922195246e-16
+ a0 = -1.385819753e+00 la0 = 1.180129697e-06 wa0 = 1.979106471e-06 pa0 = -1.041262232e-12
+ keta = -3.494008907e-01 lketa = 8.892398187e-08 wketa = 1.341030419e-07 pketa = -3.244145141e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.048960404e+00 lags = 1.356868773e-06 wags = 1.384558149e-06 pags = -9.577281044e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '3.567072202e-03+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -4.944929575e-08 wvoff = -1.042652058e-07 pvoff = 4.714129284e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.838365495e+00+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.118802841e-06 wnfactor = -2.593541421e-07 pnfactor = 1.750863609e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 9.642950748e-03 ltvoff = -5.494203926e-09 wtvoff = -5.651596932e-09 ptvoff = 2.980036997e-15
+ cit = -5.269771100e-05 lcit = 2.348656254e-11 wcit = 2.882815673e-11 pcit = -1.079902751e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.122973003e+00 leta0 = 4.855355023e-07 weta0 = 7.150999516e-07 peta0 = -2.969676022e-13
+ etab = 1.917424003e-01 letab = -6.302518720e-08 wetab = -1.297334115e-07 petab = 4.087512473e-14
+ dsub = 4.028422278e-01 ldsub = -5.619151551e-08 wdsub = -2.534656039e-08 pdsub = 1.415938250e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.152187044e+00 lpclm = -8.241274389e-07 wpclm = -9.306962907e-07 ppclm = 3.727580238e-13
+ pdiblc1 = 5.361984135e+00 lpdiblc1 = -2.069005288e-06 wpdiblc1 = -2.361848265e-06 ppdiblc1 = 9.794428754e-13
+ pdiblc2 = 3.800163548e-02 lpdiblc2 = -1.486084558e-08 wpdiblc2 = -2.242217511e-08 ppdiblc2 = 9.888850699e-15
+ pdiblcb = -0.025
+ drout = 2.120261878e+00 ldrout = -3.129641707e-07 wdrout = -8.318293337e-07 pdrout = 2.326774450e-13
+ pscbe1 = 2.849309470e+08 lpscbe1 = 6.629500152e+01 wpscbe1 = 8.512762513e+01 ppscbe1 = -4.904477695e-5
+ pscbe2 = 1.850816423e-08 lpscbe2 = -1.385706675e-15 wpscbe2 = -3.704993417e-15 ppscbe2 = 1.369159022e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.501794052e-04 lalpha0 = -4.377431138e-11 walpha0 = -4.465009890e-11 palpha0 = 1.287750770e-17
+ alpha1 = 0.0
+ beta0 = 7.501365372e+01 lbeta0 = -8.671659988e-06 wbeta0 = -1.089887611e-05 pbeta0 = 2.629710065e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -4.080308193e-06 lagidl = 1.741907519e-12 wagidl = 2.915180618e-12 pagidl = -1.119686368e-18
+ bgidl = 2.125787494e+09 lbgidl = -5.832467293e+01 wbgidl = -4.054366856e+02 pbgidl = 1.003616261e-4
+ cgidl = -8.429852818e+03 lcgidl = 3.516807801e-03 wcgidl = 6.717357163e-03 pcgidl = -2.549110444e-9
+ egidl = -5.893191400e-01 legidl = 4.314550783e-07 wegidl = 1.207686684e-06 pegidl = -3.507444222e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -8.102942212e-01 lkt1 = 1.258960579e-07 wkt1 = 2.225345482e-07 pkt1 = -1.134198317e-13
+ kt2 = -0.019032
+ at = 1.086983772e+05 lat = -4.684224981e-02 wat = -5.916028556e-02 pat = 2.807747153e-8
+ ute = -1.969877642e+00 lute = 2.204349868e-07 wute = 5.437974379e-07 pute = -2.004299506e-13
+ ua1 = 5.52e-10
+ ub1 = -1.660799783e-19 lub1 = -8.084906023e-25 wub1 = 9.811505820e-25 pub1 = -4.656540662e-31
+ uc1 = 1.211025194e-09 luc1 = -5.362038884e-16 wuc1 = -7.236473495e-16 puc1 = 3.018889738e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.38397e-10
+ cgso = 1.38397e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 7.0035e-12
+ cgdl = 7.0035e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 6.2308e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007229086434
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.322438612e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.3787656e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_g5v0d10v5
