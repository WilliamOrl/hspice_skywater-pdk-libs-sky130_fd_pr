* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param GAU = AGAUSS(0,1.0,1)
.param sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre = 0.0
* statistics '
*   process '
*   '
*   mismatch '
*     vary sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre dist=gauss std = 1.0
*   '
* '
.subckt  sky130_fd_pr__pfet_g5v0d10v5 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__pfet_g5v0d10v5 d g s b sky130_fd_pr__pfet_g5v0d10v5__model l = 'l' w = 'w' nf = 'nf' ad = 'ad' as = 'as' pd = 'pd' ps = 'ps' nrd = 'nrd' nrs = 'nrs' sa = 'sa' sb = 'sb' sd = 'sd'
.model sky130_fd_pr__pfet_g5v0d10v5__model.0 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.916781+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.0252804
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.704411452e-9
+ ub = -1.7524e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209856
+ a0 = 0.8967395
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1342734
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.1682+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.06764e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.622251
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.1 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.916781+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.0252804
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.704411452e-9
+ ub = -1.7524e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209856
+ a0 = 0.8967395
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1342734
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.1682+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.06764e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.622251
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.2 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.9182127628125+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.13241700247643e-8
+ k1 = 0.604152409375 lk1 = -7.07277513492185e-8
+ k2 = 0.02329948529375 lk2 = 1.56675496404078e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 297721.476875 lvsat = -0.772903590973594
+ ua = 2.44976570406837e-09 lua = 2.0140568818282e-15
+ ub = 8.85170975e-20 lub = -2.08612082340188e-24
+ uc = -5.15756313125e-11 luc = 9.17760209583907e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0202516383125 lu0 = 5.80508647685934e-9
+ a0 = 0.9165416104125 la0 = -1.56619841780065e-7
+ keta = -0.00495672689375 lketa = -2.34839323906078e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1097586887125 lags = 1.9389298025066e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.094776478466875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.24319289368811e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.349198275+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.43156060654374e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.64831926658375 lpclm = 5.78838869829003e-06 wpclm = 8.470329472543e-22 ppclm = -9.69352280335579e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00455412315405625 lpdiblc2 = -1.27602734399944e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 562123300.169375 lpscbe1 = -1806.55551118713
+ pscbe2 = -1.5317388699625e-08 lpscbe2 = 2.39795383634009e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.815322348125e-05 lalpha0 = -2.17393918220827e-10
+ alpha1 = 0.0
+ beta0 = 39.1402881918125 lbeta0 = -6.914600055593e-06 wbeta0 = -2.16840434497101e-19
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.570604105e-09 lagidl = -3.97806884747126e-15
+ bgidl = 1478354425.0 lbgidl = 1790.22373906875
+ cgidl = 932.600375 lcgidl = -0.00183969451596875
+ egidl = 1.20931880529938 legidl = -4.07967463450158e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.6304477199375 lkt1 = 6.4829907165672e-8
+ kt2 = -0.019032
+ at = 673047.845625 lat = -1.92232617300953
+ ute = -1.22055006875 lute = -1.31174856873906e-6
+ ua1 = 1.375495223e-09 lua1 = -5.29077591251275e-15
+ ub1 = -2.6104100625e-18 lub1 = -4.22820546317188e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.3 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.874172617125+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.60839769504094e-7
+ k1 = 0.602594105 lk1 = -6.463594997125e-8
+ k2 = 0.026832087675 lk2 = 1.85772378150623e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84545.075 lvsat = 0.06045625805625
+ ua = 3.31386607100375e-09 lua = -1.36392747761391e-15
+ ub = -1.45999138375e-18 lub = 3.96738595692469e-24 pub = 5.60519385729927e-45
+ uc = -5.4923007875e-11 luc = 1.04861752785344e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.020938342575 lu0 = 3.12058783868126e-9
+ a0 = 0.8237225450125 la0 = 2.06233089634885e-7
+ keta = -0.0050873285 lketa = -2.2973378061375e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.121306802125 lags = 1.48748517892844e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.064087020519875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.07540834542429e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.4583077875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.85809696828438e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.019094925 leta0 = 2.3809316444375e-7
+ etab = -0.1224012755 letab = 2.04849686248375e-7
+ dsub = 0.81474168125 ldsub = -9.95848917426563e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04876570365625 lpclm = -8.45940721620695e-7
+ pdiblc1 = 0.581562116725 lpdiblc1 = -7.48864204807207e-7
+ pdiblc2 = -0.001133342292 lpdiblc2 = 9.473450855001e-09 ppdiblc2 = -2.52435489670724e-29
+ pdiblcb = 0.165925 lpdiblcb = -7.4637355625e-07 wpdiblcb = 2.11758236813575e-22 ppdiblcb = 4.03896783473158e-28
+ drout = 0.139965 ldrout = 1.64202182375e-6
+ pscbe1 = -156170353.9325 lpscbe1 = 1001.43395611063 ppscbe1 = -1.73472347597681e-18
+ pscbe2 = 7.6074691134375e-08 lpscbe2 = -1.17479104457056e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.4063189874125e-05 lalpha0 = -8.41274543421732e-11
+ alpha1 = -9.54625e-11 lalpha1 = 3.73186778125e-16
+ beta0 = 70.183410779125 lbeta0 = -0.000128269927030044
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.70826975625e-09 lagidl = -6.06988294620315e-16
+ bgidl = 2620002425 lbgidl = -2672.76370493125
+ cgidl = 455.74720625 lcgidl = 2.44437339671877e-5
+ egidl = -1.5853225474425 legidl = 6.84527707370459e-06 wegidl = -1.6940658945086e-21 pegidl = -3.23117426778526e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.699418447125 lkt1 = 3.34453722423406e-7
+ kt2 = -0.019032
+ at = 210435.60875 lat = -0.113859286005938
+ ute = -1.7051169625 lute = 5.82544560653126e-7
+ ua1 = -4.84145456e-10 lua1 = 1.979024411868e-15 wua1 = -5.91645678915759e-31 pua1 = 2.25694915357879e-36
+ ub1 = -3.7199705125e-18 lub1 = 1.09343725990627e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.99339657525+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 6.67885725460622e-8
+ k1 = 0.5590564875 lk1 = 1.8488246240625e-8
+ k2 = 0.022879783675 lk2 = 9.40366019350625e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 178330.86925 lvsat = -0.118604269615563 wvsat = 8.88178419700125e-16
+ ua = 3.46201304285e-09 lua = -1.64677708361136e-15
+ ub = 4.300207475e-19 lub = 3.58880295335625e-25
+ uc = 5.32329505e-13 luc = -1.01635010742125e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.025667614225 lu0 = -5.90877405908125e-9
+ a0 = 1.02177378945 la0 = -1.71896248807413e-7
+ keta = 0.044301656 lketa = -1.17269296718e-07 pketa = -2.01948391736579e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.2888171909 lags = 9.31777751575825e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.15919953277725+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 7.40527294849646e-08 wvoff = -8.470329472543e-22
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.367170275+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 2.25157327456249e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.454625e-05 lcit = -8.6799278125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.27452410817075 leta0 = -2.49585003525004e-7
+ etab = -0.028844949 letab = 2.622726987825e-8
+ dsub = 0.0649191575000002 ldsub = 4.35749736043125e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0624965230850001 lpclm = 1.03709371138496e-6
+ pdiblc1 = -0.00178611264999995 lpdiblc1 = 3.64893402127013e-7
+ pdiblc2 = 0.005940118645525 lpdiblc2 = -4.03155443996861e-9
+ pdiblcb = -0.40685 lpdiblcb = 3.471971125e-7
+ drout = 1.5358306539575 ldrout = -1.02303467606836e-6
+ pscbe1 = 430963245.09 lpscbe1 = -119.550867823083
+ pscbe2 = 1.4532757728e-08 lpscbe2 = 1.98318990659996e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.165892571425e-05 lalpha0 = 1.17722494844932e-10 walpha0 = -5.25334031222881e-26 palpha0 = 6.33412779951888e-32
+ alpha1 = 1.90925e-10 lalpha1 = -1.7359855625e-16
+ beta0 = -39.87379705625 lbeta0 = 8.18567970296453e-05 wbeta0 = -8.13151629364128e-20 pbeta0 = 5.16987882845642e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.2060019275e-09 lagidl = 6.07971655742063e-15
+ bgidl = 855308900.0 lbgidl = 696.477407675
+ cgidl = 439.5176475 lcgidl = 5.54300190106251e-5
+ egidl = 3.11021319877 legidl = -2.11967454975162e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.64419398775 lkt1 = 2.29016423361688e-7
+ kt2 = -0.019032
+ at = 260819.25 lat = -0.2100542530625
+ ute = -1.211876175 lute = -3.59175412881251e-7
+ ua1 = 6.72948365e-10 lua1 = -2.3015696587625e-16
+ ub1 = -3.532040775e-18 lub1 = -2.49461125331251e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.5 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.91626453875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -3.34373164156219e-9
+ k1 = 0.590241525 lk1 = -9.86674910625021e-9
+ k2 = 0.02223217125 lk2 = 9.99250179093749e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8367.10762500006 lvsat = 0.0359352806419687
+ ua = -8.20535858874999e-10 lua = 2.24713050528209e-15
+ ub = 4.35210395e-18 lub = -3.2072738565375e-24 wub = -1.17549435082229e-38
+ uc = 6.082695725e-12 luc = -6.06302059295625e-18 puc = 5.87747175411144e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.019157397375 lu0 = 1.06406117812362e-11
+ a0 = 0.79446050875 la0 = 3.47883516690627e-8
+ keta = -0.1537600425 lketa = 6.2818302643125e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.78858180375 lags = -4.78472843096877e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0952545834049999+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.59107842682462e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.892981925+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.07143691530625e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.273125e-05 lcit = 1.61221390625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -7.166468125e-05 leta0 = 9.12029406765625e-11
+ etab = 0.0007545356125 letab = -6.86061505665625e-10
+ dsub = 1.499306975 ldsub = -8.6846738701875e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.0219019961875 lpclm = -7.44495715033484e-7
+ pdiblc1 = 0.1958620354125 lpdiblc1 = 1.85181823501184e-7
+ pdiblc2 = -0.033618504135125 lpdiblc2 = 3.19371233233374e-08 wpdiblc2 = -2.64697796016969e-23 ppdiblc2 = 2.52435489670724e-29
+ pdiblcb = -0.025
+ drout = 0.335842470275 ldrout = 6.80545799449564e-8
+ pscbe1 = -56987686.125 lpscbe1 = 324.118516384156
+ pscbe2 = 1.82815146225e-08 lpscbe2 = -3.38872530725812e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0002471576267875 lalpha0 = -1.63068955517284e-10
+ alpha1 = 0.0
+ beta0 = 67.19689401875 lbeta0 = -1.54972288302984e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.152563905e-08 lagidl = -1.4849134962125e-15
+ bgidl = 961697500.0 lbgidl = 599.743573125001
+ cgidl = 431.2572 lcgidl = 6.29408308999999e-5
+ egidl = 1.8355566512875 legidl = -9.60693083953159e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.4996649875 lkt1 = 9.7603429884375e-8
+ kt2 = -0.019032
+ at = 46822 lat = -0.0154772535
+ ute = -2.057628375 lute = 4.0982477496875e-7
+ ua1 = -5.03418250000002e-11 lua1 = 4.2749463938125e-16
+ ub1 = -4.570616875e-18 lub1 = 6.94864193593752e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.6 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.7943030625+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -8.98449086718752e-8
+ k1 = 0.5943829125 lk1 = -1.28040281906251e-8
+ k2 = 0.02652557625 lk2 = 6.9474042946875e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 61237.9886249999 lvsat = -0.00156339170728123
+ ua = -2.037867569625e-09 lua = 3.11052302113153e-15
+ ub = 2.53193054975e-18 lub = -1.91631587241019e-24 wub = 2.93873587705572e-39 pub = 1.40129846432482e-45
+ uc = 2.7825305e-12 luc = -3.722378407125e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00638258624999999 lu0 = 9.0711754021875e-9
+ a0 = 0.9390707625 la0 = -6.77764708031249e-8
+ keta = 0.01556431875 lketa = -5.72750005734375e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.6255407 lags = 9.55119101475e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '0.01132308791625+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.96794291163503e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.1799136+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -8.564432058e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0601722599225 leta0 = 4.27175501155331e-08 weta0 = -5.79026428787119e-24 peta0 = -3.4315449377114e-29
+ etab = -0.0007545356125 letab = 3.84247260665625e-10
+ dsub = 0.189319827725 ldsub = 6.06409971860438e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2216982981875 lpclm = 5.32298757773015e-7
+ pdiblc1 = 0.1763525393125 lpdiblc1 = 1.99018933610109e-7
+ pdiblc2 = 0.0267160385535 lpdiblc2 = -1.08551510785699e-8
+ pdiblcb = -0.025
+ drout = -0.738324518225 ldrout = 8.29907516538581e-7
+ pscbe1 = 432224423.35 lpscbe1 = -22.8551722609875
+ pscbe2 = 1.054562873625e-08 lpscbe2 = 2.09795175756469e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.00012163830041875 lalpha0 = 9.84995558537484e-11 walpha0 = 2.06795153138257e-25 palpha0 = 9.86076131526265e-32
+ alpha1 = 0.0
+ beta0 = 26.4659450525 lbeta0 = 1.33911967240144e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.84437134625e-08 lagidl = -6.39155777327812e-15 wagidl = 1.0097419586829e-28
+ bgidl = 2062179625 lbgidl = -180.77337403125
+ cgidl = 1258.4125 lcgidl = -0.000523719065625
+ egidl = -0.2467454455 legidl = 5.16179678193375e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.0943169337500003 lkt1 = -3.23678247762188e-7
+ kt2 = -0.019032
+ at = 42823.75 lat = -0.0126414946875
+ ute = -1.613478125 lute = 9.48112101562502e-8
+ ua1 = 5.534185e-10 lua1 = -7.22371124999967e-19
+ ub1 = -4.333641125e-18 lub1 = 5.26789142906249e-25
+ uc1 = -2.8159131e-10 luc1 = 1.222685366175e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.7 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 2.0e-05 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.842322719999999+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -6.53908980900007e-8
+ k1 = 0.451376 lk1 = 6.00222420000003e-8
+ k2 = 0.0478496225 lk2 = -3.91186625812501e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 38528.5017499999 lvsat = 0.0100014144838125
+ ua = 1.188723724875e-08 lua = -3.98083660762594e-15
+ ub = -8.64438477450001e-18 lub = 3.77522270646413e-24 pub = 1.12103877145985e-44
+ uc = -1.43920875e-12 luc = -1.5724576940625e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03876347225 lu0 = -7.41879079331252e-9
+ a0 = 0.177126449999999 la0 = 3.202436703375e-7
+ keta = -0.1420657375 lketa = 2.29981055718751e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.123592234725+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 9.02619893870631e-9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.440028875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -4.79656909593749e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.04625e-05 lcit = -1.0420528125e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.20687682 leta0 = 1.17426847335e-07 peta0 = -2.01948391736579e-28
+ etab = 0.01575735275 letab = -8.02443188793751e-9
+ dsub = 0.42597171955 ldsub = -5.98739787258376e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.98195066125 lpclm = 1.45140241883437e-7
+ pdiblc1 = 1.6849454761 lpdiblc1 = -5.69232019448926e-7
+ pdiblc2 = 0.00785230350750001 lpdiblc2 = -1.24879400639438e-9
+ pdiblcb = -0.025
+ drout = 0.85752593545 ldrout = 1.72206730045875e-8
+ pscbe1 = 488447117 lpscbe1 = -51.4865790022501
+ pscbe2 = 1.539618939e-08 lpscbe2 = -3.72196255357505e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.19739062200001e-05 lalpha0 = 5.28379631080351e-11
+ alpha1 = 0.0
+ beta0 = 44.8934311525 lbeta0 = 4.00699942758938e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -4.9973592500001e-10 lagidl = 3.25539382730626e-15
+ bgidl = 2086574750 lbgidl = -193.1965914375
+ cgidl = -2413.755 lcgidl = 0.00134633223375 pcgidl = -1.65436122510606e-24
+ egidl = 1.1826331595 legidl = -2.11731376402875e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.943332292500001 lkt1 = 2.04744620705625e-7
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.65197825 lute = 1.144173988125e-7
+ ua1 = 5.52e-10
+ ub1 = -7.96137600000001e-18 lub1 = 2.374213128e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.8 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.916781+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.0252804
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.704411452e-9
+ ub = -1.7524e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209856
+ a0 = 0.8967395
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1342734
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.1682+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.06764e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.622251
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.9 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.916781+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.0252804
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.704411452e-9
+ ub = -1.7524e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209856
+ a0 = 0.8967395
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1342734
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.1682+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.06764e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.622251
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.10 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.9182127628125+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.13241700247643e-8
+ k1 = 0.604152409375001 lk1 = -7.07277513492185e-8
+ k2 = 0.02329948529375 lk2 = 1.56675496404078e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 297721.476875 lvsat = -0.772903590973594
+ ua = 2.44976570406837e-09 lua = 2.01405688182821e-15
+ ub = 8.85170974999998e-20 lub = -2.08612082340187e-24 pub = 1.12103877145985e-44
+ uc = -5.15756313125e-11 luc = 9.17760209583907e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0202516383125 lu0 = 5.80508647685937e-9
+ a0 = 0.9165416104125 la0 = -1.56619841780065e-7
+ keta = -0.00495672689375 lketa = -2.34839323906078e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1097586887125 lags = 1.93892980250659e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0947764784668749+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.24319289368814e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.349198275+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.43156060654375e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.64831926658375 lpclm = 5.78838869829003e-06 wpclm = 3.3881317890172e-21 ppclm = -6.46234853557053e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00455412315405625 lpdiblc2 = -1.27602734399944e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 562123300.169375 lpscbe1 = -1806.55551118713
+ pscbe2 = -1.5317388699625e-08 lpscbe2 = 2.39795383634009e-13 ppscbe2 = 7.70371977754894e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.815322348125e-05 lalpha0 = -2.17393918220827e-10
+ alpha1 = 0.0
+ beta0 = 39.1402881918125 lbeta0 = -6.91460005559311e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.570604105e-09 lagidl = -3.97806884747124e-15
+ bgidl = 1478354425.0 lbgidl = 1790.22373906875
+ cgidl = 932.600375 lcgidl = -0.00183969451596875
+ egidl = 1.20931880529937 legidl = -4.07967463450158e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.630447719937501 lkt1 = 6.4829907165672e-8
+ kt2 = -0.019032
+ at = 673047.845625 lat = -1.92232617300953
+ ute = -1.22055006875 lute = -1.31174856873907e-6
+ ua1 = 1.375495223e-09 lua1 = -5.29077591251275e-15
+ ub1 = -2.6104100625e-18 lub1 = -4.22820546317187e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.11 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.874172617125+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.60839769504093e-7
+ k1 = 0.602594105 lk1 = -6.46359499712504e-8
+ k2 = 0.026832087675 lk2 = 1.85772378150626e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84545.075 lvsat = 0.0604562580562502
+ ua = 3.31386607100375e-09 lua = -1.36392747761392e-15
+ ub = -1.45999138375e-18 lub = 3.96738595692469e-24 pub = 1.12103877145985e-44
+ uc = -5.4923007875e-11 luc = 1.04861752785344e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.020938342575 lu0 = 3.12058783868126e-9
+ a0 = 0.8237225450125 la0 = 2.06233089634883e-7
+ keta = -0.0050873285 lketa = -2.2973378061375e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.121306802125 lags = 1.48748517892844e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0640870205198749+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.07540834542429e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.4583077875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.85809696828437e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.019094925 leta0 = 2.3809316444375e-7
+ etab = -0.1224012755 letab = 2.04849686248375e-7
+ dsub = 0.81474168125 ldsub = -9.95848917426562e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04876570365625 lpclm = -8.45940721620696e-07 wpclm = -1.35525271560688e-20
+ pdiblc1 = 0.581562116725 lpdiblc1 = -7.48864204807207e-7
+ pdiblc2 = -0.001133342292 lpdiblc2 = 9.47345085500101e-9
+ pdiblcb = 0.165925 lpdiblcb = -7.4637355625e-07 wpdiblcb = -8.470329472543e-22 ppdiblcb = 2.42338070083895e-27
+ drout = 0.139965 ldrout = 1.64202182375e-6
+ pscbe1 = -156170353.9325 lpscbe1 = 1001.43395611063
+ pscbe2 = 7.6074691134375e-08 lpscbe2 = -1.17479104457055e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.4063189874125e-05 lalpha0 = -8.41274543421732e-11
+ alpha1 = -9.54625e-11 lalpha1 = 3.73186778125e-16
+ beta0 = 70.183410779125 lbeta0 = -0.000128269927030044
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.70826975625e-09 lagidl = -6.06988294620309e-16
+ bgidl = 2620002425.0 lbgidl = -2672.76370493125
+ cgidl = 455.74720625 lcgidl = 2.44437339671881e-5
+ egidl = -1.5853225474425 legidl = 6.84527707370459e-06 wegidl = 3.3881317890172e-21 pegidl = 1.93870456067116e-26
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.699418447125001 lkt1 = 3.34453722423406e-7
+ kt2 = -0.019032
+ at = 210435.60875 lat = -0.113859286005937
+ ute = -1.7051169625 lute = 5.82544560653127e-7
+ ua1 = -4.84145456e-10 lua1 = 1.979024411868e-15 wua1 = -1.57772181044202e-30 pua1 = -9.02779661431517e-36
+ ub1 = -3.7199705125e-18 lub1 = 1.09343725990636e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.12 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.984047538342441+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 4.89389238303069e-08 wvth0 = -1.86751181898939e-07 pvth0 = 3.56554694040543e-13
+ k1 = 0.5590564875 lk1 = 1.8488246240625e-8
+ k2 = 0.0232555969850038 lk2 = 8.68613863138151e-09 wk2 = -7.50703848006211e-09 pk2 = 1.43328132180586e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 178330.86925 lvsat = -0.118604269615563
+ ua = 3.45991826490661e-09 lua = -1.64277762882294e-15 wua = 4.18441236902234e-17 pua = -7.989089315553e-23
+ ub = 3.46306971054226e-19 lub = 5.18710823014719e-25 wub = 1.67222002084863e-24 pub = -3.19268607480524e-30
+ uc = 5.32329505e-13 luc = -1.01635010742125e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0251605385849804 lu0 = -4.94063989337381e-09 wu0 = 1.01290620651274e-08 pu0 = -1.93389117478444e-14
+ a0 = 1.02109296823622 la0 = -1.70596390905012e-07 wa0 = 1.35997073914275e-08 pa0 = -2.59652413370807e-14
+ keta = 0.044301656 lketa = -1.17269296718e-07 pketa = 4.03896783473158e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.284887490854091 lags = 9.24274971763173e-07 wags = -7.84975110632591e-08 pags = 1.49871372997517e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.15919953277725+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 7.40527294849646e-08 wvoff = -1.6940658945086e-21
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.99590485070422+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 9.33995838792968e-07 wnfactor = 7.41619243468743e-06 pnfactor = -1.41593654059271e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.454625e-05 lcit = -8.67992781250001e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.274560812604027 leta0 = -2.49655081464239e-07 weta0 = -7.3318742488618e-10 peta0 = 1.39983809096307e-15
+ etab = -0.028844949 letab = 2.622726987825e-8
+ dsub = 0.0649191575000003 ldsub = 4.35749736043125e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0624965230849996 lpclm = 1.03709371138496e-6
+ pdiblc1 = -0.00178611265000006 lpdiblc1 = 3.64893402127013e-7
+ pdiblc2 = 0.005940118645525 lpdiblc2 = -4.03155443996861e-09 ppdiblc2 = 5.04870979341448e-29
+ pdiblcb = -0.40685 lpdiblcb = 3.471971125e-7
+ drout = 1.5358306539575 ldrout = -1.02303467606836e-6
+ pscbe1 = 430963245.09 lpscbe1 = -119.550867823083
+ pscbe2 = 1.4532757728e-08 lpscbe2 = 1.98318990660185e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.165892571425e-05 lalpha0 = 1.17722494844932e-10 walpha0 = -5.11797178089288e-26 palpha0 = 3.15079129636214e-31
+ alpha1 = 1.90925e-10 lalpha1 = -1.7359855625e-16
+ beta0 = -39.87379705625 lbeta0 = 8.18567970296453e-05 wbeta0 = -1.0842021724855e-19 pbeta0 = -5.16987882845642e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -4.47480514352114e-09 lagidl = 2.07442974577677e-14 wagidl = 1.53427546883601e-13 pagidl = -2.92931543887515e-19
+ bgidl = 1039402956.20476 lbgidl = 344.995830866063 wbgidl = -3677.36087863913 pbgidl = 0.00702100125754179
+ cgidl = 78.7368698963523 lcgidl = 0.000744250718650389 wcgidl = 0.00720675694085968 pcgidl = -1.37595006893363e-8
+ egidl = 3.11021319877 legidl = -2.11967454975162e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.357323161113766 lkt1 = -3.18691702393541e-07 wkt1 = -5.73037270644744e-06 pkt1 = 1.09407140897848e-11
+ kt2 = -0.019032
+ at = 266265.8197102 lat = -0.2204531162817 wat = -0.108797659131334 pat = 2.07721930696504e-7
+ ute = -1.211876175 lute = -3.5917541288125e-7
+ ua1 = 6.72948365e-10 lua1 = -2.3015696587625e-16
+ ub1 = -3.532040775e-18 lub1 = -2.49461125331251e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.13 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.96300972328779+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 2.98102904918669e-08 wvth0 = 9.33755909494666e-07 pvth0 = -6.62266378809097e-13
+ k1 = 0.590241525000001 lk1 = -9.86674910625021e-9
+ k2 = 0.020353104699981 lk2 = 1.13252297415385e-08 wk2 = 3.75351924003118e-08 pk2 = -2.66218352099206e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8367.10762500006 lvsat = 0.0359352806419687
+ ua = -8.1006196915804e-10 lua = 2.23970189900034e-15 wua = -2.09220618451016e-16 pua = 1.48389723636375e-22
+ ub = 4.77067283222887e-18 lub = -3.50414383625833e-24 wub = -8.36110010424311e-24 pub = 5.93011024893446e-30
+ uc = 6.08269572499999e-12 luc = -6.06302059295625e-18 puc = -2.35098870164458e-38
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0216927755750981 lu0 = -1.78757637663835e-09 wu0 = -5.06453103256378e-08 pu0 = 3.59201863484578e-14
+ a0 = 0.797864614818877 la0 = 3.23739894397137e-08 wa0 = -6.79985369571106e-08 pa0 = 4.82279623368387e-14
+ keta = -0.1537600425 lketa = 6.28183026431248e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.768933303520454 lags = -3.39115855218822e-08 wags = 3.92487555316262e-07 pags = -2.78371798608083e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0952545834049998+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.59107842682461e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '7.74930904647891+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -3.38803692621516e-06 wnfactor = -3.70809621734374e-05 pnfactor = 2.62996724215105e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.273125e-05 lcit = 1.61221390625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.000255186847635189 leta0 = 2.21366037185258e-10 weta0 = 3.66593712443036e-09 peta0 = -2.60006590550223e-15
+ etab = 0.0007545356125 letab = -6.86061505665625e-10
+ dsub = 1.499306975 ldsub = -8.68467387018751e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.0219019961875 lpclm = -7.44495715033487e-7
+ pdiblc1 = 0.1958620354125 lpdiblc1 = 1.85181823501184e-7
+ pdiblc2 = -0.033618504135125 lpdiblc2 = 3.19371233233374e-08 wpdiblc2 = 1.05879118406788e-22 ppdiblc2 = 1.51461293802434e-28
+ pdiblcb = -0.025
+ drout = 0.335842470275 ldrout = 6.80545799449566e-8
+ pscbe1 = -56987686.125 lpscbe1 = 324.118516384157
+ pscbe2 = 1.82815146225e-08 lpscbe2 = -3.38872530725811e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0002471576267875 lalpha0 = -1.63068955517284e-10
+ alpha1 = 0.0
+ beta0 = 67.1968940187498 lbeta0 = -1.54972288302985e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.99296744051057e-08 lagidl = -2.87229755718212e-14 wagidl = -7.67137734418005e-13 pagidl = 5.4409243813597e-19
+ bgidl = 41227218.9761963 lbgidl = 1252.58711994113 wbgidl = 18386.8043931957 pbgidl = -0.0130408410158741
+ cgidl = 2235.16108801824 lcgidl = -0.00121647800167694 wcgidl = -0.0360337847042984 pcgidl = 2.55569618015237e-8
+ egidl = 1.8355566512875 legidl = -9.60693083953159e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.93401912068117 lkt1 = 1.11491909884312e-06 wkt1 = 2.86518635322373e-05 pkt1 = -2.03213342102393e-11
+ kt2 = -0.019032
+ at = 19589.1514489999 lat = 0.00383764433479683 wat = 0.54398829565668 pat = -3.85823698694499e-7
+ ute = -2.057628375 lute = 4.09824774968749e-7
+ ua1 = -5.03418250000006e-11 lua1 = 4.2749463938125e-16
+ ub1 = -4.57061687500001e-18 lub1 = 6.94864193593755e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.14 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.794303062499999+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -8.98449086718761e-8
+ k1 = 0.594382912500001 lk1 = -1.28040281906247e-8
+ k2 = 0.0265255762500001 lk2 = 6.94740429468753e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 61237.988625 lvsat = -0.00156339170728126
+ ua = -2.037867569625e-09 lua = 3.11052302113153e-15
+ ub = 2.53193054975e-18 lub = -1.91631587241019e-24 wub = -5.87747175411144e-39 pub = 8.4077907859489e-45
+ uc = 2.78253049999999e-12 luc = -3.722378407125e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00638258625000004 lu0 = 9.07117540218748e-9
+ a0 = 0.9390707625 la0 = -6.77764708031244e-8
+ keta = 0.01556431875 lketa = -5.72750005734375e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.6255407 lags = 9.55119101474999e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '0.0113230879162498+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.96794291163503e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.17991360000001+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -8.56443205799999e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0601722599225 leta0 = 4.27175501155331e-08 weta0 = -9.76073122812573e-23 peta0 = 4.25984888819346e-29
+ etab = -0.0007545356125 letab = 3.84247260665625e-10
+ dsub = 0.189319827725 ldsub = 6.06409971860439e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2216982981875 lpclm = 5.32298757773016e-7
+ pdiblc1 = 0.1763525393125 lpdiblc1 = 1.99018933610109e-7
+ pdiblc2 = 0.0267160385535 lpdiblc2 = -1.08551510785699e-8
+ pdiblcb = -0.025
+ drout = -0.738324518224999 ldrout = 8.29907516538581e-7
+ pscbe1 = 432224423.350001 lpscbe1 = -22.8551722609877
+ pscbe2 = 1.054562873625e-08 lpscbe2 = 2.09795175756468e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.00012163830041875 lalpha0 = 9.84995558537484e-11 walpha0 = 4.13590306276514e-25 palpha0 = 3.94430452610506e-31
+ alpha1 = 0.0
+ beta0 = 26.4659450525 lbeta0 = 1.33911967240144e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.84437134625e-08 lagidl = -6.39155777327813e-15
+ bgidl = 2062179625 lbgidl = -180.773374031251
+ cgidl = 1258.4125 lcgidl = -0.000523719065625 pcgidl = -6.61744490042422e-24
+ egidl = -0.2467454455 legidl = 5.16179678193375e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.0943169337500001 lkt1 = -3.23678247762188e-7
+ kt2 = -0.019032
+ at = 42823.75 lat = -0.0126414946875
+ ute = -1.613478125 lute = 9.48112101562498e-8
+ ua1 = 5.53418500000001e-10 lua1 = -7.22371125000165e-19
+ ub1 = -4.333641125e-18 lub1 = 5.26789142906249e-25
+ uc1 = -2.8159131e-10 luc1 = 1.222685366175e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.15 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-05 wmax = 2.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.765544801901044+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.04490052881893e-07 wvth0 = -1.53367315697809e-06 pvth0 = 7.81023055191092e-13
+ k1 = 0.451376 lk1 = 6.00222420000003e-8
+ k2 = 0.0466361396474511 lk2 = -3.2939001154645e-09 wk2 = 2.42398611930178e-08 pk2 = -1.23441493125445e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 44207.3563518783 lvsat = 0.00710945777780603 wvsat = -0.113437653441672 pvsat = 5.7768125015172e-8
+ ua = 1.1878881254857e-08 lua = -3.97658131773591e-15 wua = 1.66914704786938e-16 pua = -8.50013134126814e-23
+ ub = -8.54938990472976e-18 lub = 3.72684656903363e-24 wub = -1.89756489137272e-24 pub = 9.66334920931517e-31
+ uc = -1.43920874999999e-12 luc = -1.5724576940625e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0361305821820452 lu0 = -6.07799152620649e-09 wu0 = 5.25931533763674e-08 pu0 = -2.67830633569153e-14
+ a0 = 0.177126449999999 la0 = 3.202436703375e-7
+ keta = -0.1420657375 lketa = 2.29981055718751e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.123592234725+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 9.02619893870626e-9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.07945646619626+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.31453541041044e-06 wnfactor = -3.27482973188509e-05 pnfactor = 1.66770704096248e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.04625e-05 lcit = -1.0420528125e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.344257787791609 leta0 = 1.87388105182877e-07 weta0 = 2.74424610354902e-06 peta0 = -1.39750732823234e-12
+ etab = 0.01575735275 letab = -8.02443188793751e-9
+ dsub = 0.425971719550001 ldsub = -5.98739787258377e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.98195066125 lpclm = 1.45140241883437e-7
+ pdiblc1 = 1.6849454761 lpdiblc1 = -5.69232019448926e-7
+ pdiblc2 = 0.00785230350750001 lpdiblc2 = -1.24879400639438e-9
+ pdiblcb = -0.025
+ drout = 0.857525935449999 ldrout = 1.72206730045871e-8
+ pscbe1 = 488447117.0 lpscbe1 = -51.4865790022504
+ pscbe2 = 1.53961893900001e-08 lpscbe2 = -3.72196255357492e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.19739062200001e-05 lalpha0 = 5.28379631080351e-11
+ alpha1 = 0.0
+ beta0 = 44.8934311525002 lbeta0 = 4.00699942758944e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.13814109846004e-09 lagidl = 6.12675166189078e-15 wagidl = 1.12629658068571e-13 pagidl = -5.735665337142e-20
+ bgidl = 2147861762.755 lbgidl = -224.407002682983 wbgidl = -1224.23541378882 pbgidl = 0.000623441884471942
+ cgidl = -9269.56539482535 lcgidl = 0.00483765367731481 wcgidl = 0.136947870328072 pcgidl = -6.97407029645709e-8
+ egidl = 1.1826331595 legidl = -2.11731376402875e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.603066797684239 lkt1 = 3.14644174706984e-08 wkt1 = -6.79695501735553e-06 pkt1 = 3.46134934258829e-12
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.65197825 lute = 1.14417398812498e-7
+ ua1 = 5.52e-10
+ ub1 = -7.961376e-18 lub1 = 2.374213128e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.16 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.916781+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.0252804
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.704411452e-9
+ ub = -1.7524e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209856
+ a0 = 0.8967395
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1342734
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.1682+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.06764e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.622251
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.17 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.916781+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.0252804
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.704411452e-9
+ ub = -1.7524e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209856
+ a0 = 0.8967395
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1342734
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.1682+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.06764e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.622251
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.18 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.918212762812499+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.13241700247643e-8
+ k1 = 0.604152409375 lk1 = -7.07277513492202e-8
+ k2 = 0.02329948529375 lk2 = 1.56675496404079e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 297721.476875 lvsat = -0.772903590973594 wvsat = 1.77635683940025e-15
+ ua = 2.44976570406837e-09 lua = 2.01405688182821e-15
+ ub = 8.85170975000002e-20 lub = -2.08612082340188e-24 pub = -5.60519385729927e-45
+ uc = -5.15756313125e-11 luc = 9.17760209583907e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0202516383125 lu0 = 5.80508647685926e-9
+ a0 = 0.9165416104125 la0 = -1.56619841780065e-7
+ keta = -0.00495672689374999 lketa = -2.34839323906078e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1097586887125 lags = 1.93892980250659e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.094776478466875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.2431928936881e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.349198275+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.43156060654374e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.64831926658375 lpclm = 5.78838869829003e-06 ppclm = -3.23117426778526e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00455412315405625 lpdiblc2 = -1.27602734399944e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 562123300.169375 lpscbe1 = -1806.55551118713
+ pscbe2 = -1.5317388699625e-08 lpscbe2 = 2.39795383634009e-13 ppscbe2 = 3.85185988877447e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.815322348125e-05 lalpha0 = -2.17393918220827e-10
+ alpha1 = 0.0
+ beta0 = 39.1402881918125 lbeta0 = -6.914600055593e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.570604105e-09 lagidl = -3.97806884747127e-15
+ bgidl = 1478354425.0 lbgidl = 1790.22373906875
+ cgidl = 932.600375 lcgidl = -0.00183969451596875
+ egidl = 1.20931880529938 legidl = -4.07967463450159e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.6304477199375 lkt1 = 6.48299071656703e-8
+ kt2 = -0.019032
+ at = 673047.845625 lat = -1.92232617300953
+ ute = -1.22055006875 lute = -1.31174856873906e-6
+ ua1 = 1.375495223e-09 lua1 = -5.29077591251275e-15
+ ub1 = -2.6104100625e-18 lub1 = -4.22820546317189e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.19 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.874172617125+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.60839769504095e-7
+ k1 = 0.602594105 lk1 = -6.46359499712504e-8
+ k2 = 0.026832087675 lk2 = 1.85772378150631e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84545.075 lvsat = 0.06045625805625
+ ua = 3.31386607100375e-09 lua = -1.36392747761391e-15
+ ub = -1.45999138375e-18 lub = 3.96738595692469e-24 pub = -5.60519385729927e-45
+ uc = -5.4923007875e-11 luc = 1.04861752785344e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.020938342575 lu0 = 3.12058783868126e-9
+ a0 = 0.8237225450125 la0 = 2.06233089634885e-7
+ keta = -0.00508732850000001 lketa = -2.2973378061375e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.121306802125 lags = 1.48748517892844e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.064087020519875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.07540834542429e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.4583077875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.85809696828438e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.019094925 leta0 = 2.3809316444375e-7
+ etab = -0.1224012755 letab = 2.04849686248375e-7
+ dsub = 0.81474168125 ldsub = -9.95848917426563e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04876570365625 lpclm = -8.45940721620696e-7
+ pdiblc1 = 0.581562116725 lpdiblc1 = -7.48864204807206e-7
+ pdiblc2 = -0.001133342292 lpdiblc2 = 9.473450855001e-9
+ pdiblcb = 0.165925 lpdiblcb = -7.4637355625e-07 wpdiblcb = 2.11758236813575e-22
+ drout = 0.139965 ldrout = 1.64202182375e-6
+ pscbe1 = -156170353.9325 lpscbe1 = 1001.43395611063 ppscbe1 = 1.73472347597681e-18
+ pscbe2 = 7.6074691134375e-08 lpscbe2 = -1.17479104457056e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.4063189874125e-05 lalpha0 = -8.41274543421731e-11
+ alpha1 = -9.54625e-11 lalpha1 = 3.73186778125e-16
+ beta0 = 70.183410779125 lbeta0 = -0.000128269927030044
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.70826975624999e-09 lagidl = -6.06988294620309e-16
+ bgidl = 2620002425.0 lbgidl = -2672.76370493125
+ cgidl = 455.74720625 lcgidl = 2.44437339671872e-5
+ egidl = -1.5853225474425 legidl = 6.84527707370459e-06 wegidl = 1.6940658945086e-21 pegidl = -6.46234853557053e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.699418447125 lkt1 = 3.34453722423407e-7
+ kt2 = -0.019032
+ at = 210435.60875 lat = -0.113859286005938
+ ute = -1.7051169625 lute = 5.82544560653127e-7
+ ua1 = -4.84145456e-10 lua1 = 1.979024411868e-15 wua1 = 9.86076131526265e-31 pua1 = 4.89005649942072e-36
+ ub1 = -3.7199705125e-18 lub1 = 1.09343725990624e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.20 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.986783919467533+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 5.41633594933882e-08 wvth0 = -1.45772654124708e-07 pvth0 = 2.78316439887601e-13
+ k1 = 0.5590564875 lk1 = 1.84882462406254e-8
+ k2 = 0.0221266511151354 lk2 = 1.08415785334277e-08 wk2 = 9.3994294310752e-09 pk2 = -1.79458606412801e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 178330.86925 lvsat = -0.118604269615563
+ ua = 3.46147924147713e-09 lua = -1.64575792334021e-15 wua = 1.84678033511199e-17 pua = -3.52596535481094e-23
+ ub = 2.70254765694252e-19 lub = 6.6391349609825e-25 wub = 2.81113571539783e-24 pub = -5.36716086462331e-30
+ uc = 5.32329505e-13 luc = -1.01635010742125e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0243002476492448 lu0 = -3.29812942432061e-09 wu0 = 2.3012302517525e-08 pu0 = -4.39362385815849e-14
+ a0 = 1.00778995289515 la0 = -1.45197608865059e-07 wa0 = 2.12818295268911e-07 pa0 = -4.06323330242158e-13
+ keta = 0.044301656 lketa = -1.17269296718e-07 pketa = -1.0097419586829e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.311291769269596 lags = 9.74687340327977e-07 wags = 3.16918334517115e-07 pags = -6.05076330176797e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.15919953277725+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 7.40527294849647e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.32454550675617+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 3.06538666225787e-07 wnfactor = 2.49465203657696e-06 pnfactor = -4.76291440083457e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.454625e-05 lcit = -8.6799278125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.27451185329925 leta0 = -2.49561605911593e-7
+ etab = -0.028844949 letab = 2.622726987825e-8
+ dsub = 0.0649191575000001 ldsub = 4.35749736043125e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0625191985206888 lpclm = 1.03705041830938e-06 wpclm = -3.39574762684141e-10 ppclm = 6.48333115648567e-16
+ pdiblc1 = -0.00178611264999984 lpdiblc1 = 3.64893402127012e-7
+ pdiblc2 = 0.005940118645525 lpdiblc2 = -4.03155443996861e-9
+ pdiblcb = -0.40685 lpdiblcb = 3.471971125e-7
+ drout = 1.5358306539575 ldrout = -1.02303467606836e-6
+ pscbe1 = 430963245.09 lpscbe1 = -119.550867823083
+ pscbe2 = 1.4532757728e-08 lpscbe2 = 1.98318990659932e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.165892571425e-05 lalpha0 = 1.17722494844932e-10 walpha0 = 9.34003423172626e-26 palpha0 = 1.14201627171087e-31
+ alpha1 = 1.90925e-10 lalpha1 = -1.7359855625e-16
+ beta0 = -39.87379705625 lbeta0 = 8.18567970296453e-05 wbeta0 = -2.71050543121376e-20 pbeta0 = -7.75481824268463e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.29376702483197e-09 lagidl = 5.91215104533957e-15 wagidl = 3.70897138793261e-14 pagidl = -7.08135362241033e-20
+ bgidl = 793843600.0 lbgidl = 813.830031700001
+ cgidl = 559.9750875 lcgidl = -0.000174553348309375
+ egidl = 3.11021319877 legidl = -2.11967454975162e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.740627435297836 lkt1 = 4.13131983092393e-07 wkt1 = 9.77975316527818e-09 pkt1 = -1.86719937308106e-14
+ kt2 = -0.019032
+ at = 255735.48726082 lat = -0.200348079052721 wat = 0.0488987658264026 pat = -9.33599686540571e-8
+ ute = -0.94684568266989 lute = -8.65184880362511e-07 wute = -3.96894982624298e-06 pute = 7.57771745575441e-12
+ ua1 = 9.13453106089158e-10 lua1 = -6.89340642800725e-16 wua1 = -3.60166576292467e-15 pua1 = 6.87648035786392e-21
+ ub1 = -3.14111626372595e-18 lub1 = -9.95833748481232e-25 wub1 = -5.85426890866095e-24 pub1 = 1.11772629138609e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.21 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.949327817662331+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 2.01063989270087e-08 wvth0 = 7.28863270623548e-07 pvth0 = -5.16946274689734e-13
+ k1 = 0.590241525 lk1 = -9.86674910625021e-9
+ k2 = 0.025997834049323 lk2 = 7.32170545051759e-09 wk2 = -4.69971471553751e-08 pk2 = 3.33327266199498e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8367.10762499995 lvsat = 0.0359352806419688
+ ua = -8.17866852010644e-10 lua = 2.24523751216355e-15 wua = -9.23390167555488e-17 pua = 6.54914476338717e-23
+ ub = 5.15093385902874e-18 lub = -3.77384396951613e-24 wub = -1.40556785769891e-23 pub = 9.96899003072955e-30
+ uc = 6.082695725e-12 luc = -6.06302059295625e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.025994230253776 lu0 = -4.83838310749067e-09 wu0 = -1.15061512587626e-07 pu0 = 8.16073778027737e-14
+ a0 = 0.864379691524267 la0 = -1.48018287135877e-08 wa0 = -1.06409147634454e-06 pa0 = 7.54706879597368e-13
+ keta = -0.1537600425 lketa = 6.2818302643125e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.900954695597985 lags = -1.27547757852869e-07 wags = -1.58459167258558e-06 pags = 1.12387164378132e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0952545834049999+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.59107842682462e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '6.10610576621917+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.22259499969094e-06 wnfactor = -1.24732601828848e-05 pnfactor = 8.84665978471103e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.273125e-05 lcit = 1.61221390625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.039032375e-05 leta0 = 4.77441026196875e-11
+ etab = 0.0007545356125 letab = -6.86061505665625e-10
+ dsub = 1.499306975 ldsub = -8.6846738701875e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.02178861900905 lpclm = -7.44415302269674e-07 wpclm = 1.69787381341393e-09 ppclm = -1.20421700215833e-15
+ pdiblc1 = 0.1958620354125 lpdiblc1 = 1.85181823501185e-7
+ pdiblc2 = -0.033618504135125 lpdiblc2 = 3.19371233233374e-08 wpdiblc2 = -2.64697796016969e-23 ppdiblc2 = -2.52435489670724e-29
+ pdiblcb = -0.025
+ drout = 0.335842470275001 ldrout = 6.80545799449566e-8
+ pscbe1 = -56987686.125 lpscbe1 = 324.118516384156
+ pscbe2 = 1.82815146225e-08 lpscbe2 = -3.38872530725811e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0002471576267875 lalpha0 = -1.63068955517284e-10
+ alpha1 = 0.0
+ beta0 = 67.1968940187501 lbeta0 = -1.54972288302985e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.10868135633401e-08 lagidl = -1.173676519799e-15 wagidl = -1.8544856939663e-13 pagidl = 1.3152939784456e-19
+ bgidl = 1269024000.0 lbgidl = 381.772252999999
+ cgidl = -171.03 lcgidl = 0.000490113027500001
+ egidl = 1.8355566512875 legidl = -9.6069308395316e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.0174977497608206 lkt1 = -2.44373683482138e-07 wkt1 = -4.88987658264011e-08 pkt1 = 3.4681449662373e-14
+ kt2 = -0.019032
+ at = 72240.8136959 lat = -0.0335055471138171 wat = -0.24449382913201 pat = 1.73407248311879e-7
+ ute = -3.38278083665055 lute = 1.3496891583944e-06 wute = 1.98447491312149e-05 pute = -1.40748883213141e-11
+ ua1 = -1.25286553044579e-09 lua1 = 1.28038457746868e-15 wua1 = 1.80083288146233e-14 pua1 = -1.27724072117716e-20
+ ub1 = -6.52523943137025e-18 lub1 = 2.08118024169935e-24 wub1 = 2.92713445433046e-23 pub1 = -2.07607011173388e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.22 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.794303062499999+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -8.98449086718752e-8
+ k1 = 0.5943829125 lk1 = -1.28040281906251e-8
+ k2 = 0.02652557625 lk2 = 6.94740429468753e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 61237.988625 lvsat = -0.00156339170728126
+ ua = -2.037867569625e-09 lua = 3.11052302113153e-15
+ ub = 2.53193054975e-18 lub = -1.91631587241019e-24 pub = -4.20389539297445e-45
+ uc = 2.7825305e-12 luc = -3.722378407125e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00638258625000002 lu0 = 9.07117540218748e-9
+ a0 = 0.9390707625 la0 = -6.77764708031244e-8
+ keta = 0.0155643187500001 lketa = -5.72750005734375e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.625540699999999 lags = 9.55119101474999e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '0.0113230879162499+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.96794291163503e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.1799136+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -8.564432058e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0601722599225 leta0 = 4.27175501155331e-08 weta0 = -1.05051937794235e-22 peta0 = -7.80972296168802e-29
+ etab = -0.0007545356125 letab = 3.84247260665625e-10
+ dsub = 0.189319827725 ldsub = 6.06409971860436e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2216982981875 lpclm = 5.32298757773015e-7
+ pdiblc1 = 0.176352539312501 lpdiblc1 = 1.99018933610109e-7
+ pdiblc2 = 0.0267160385535 lpdiblc2 = -1.08551510785699e-8
+ pdiblcb = -0.025
+ drout = -0.738324518224998 ldrout = 8.29907516538581e-7
+ pscbe1 = 432224423.35 lpscbe1 = -22.8551722609877
+ pscbe2 = 1.054562873625e-08 lpscbe2 = 2.09795175756468e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.00012163830041875 lalpha0 = 9.84995558537484e-11 walpha0 = -2.06795153138257e-25 palpha0 = 1.97215226305253e-31
+ alpha1 = 0.0
+ beta0 = 26.4659450525 lbeta0 = 1.33911967240144e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.84437134625e-08 lagidl = -6.39155777327813e-15
+ bgidl = 2062179625.0 lbgidl = -180.773374031251
+ cgidl = 1258.4125 lcgidl = -0.000523719065625
+ egidl = -0.246745445499999 legidl = 5.16179678193375e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.0943169337500001 lkt1 = -3.23678247762187e-7
+ kt2 = -0.019032
+ at = 42823.75 lat = -0.0126414946875
+ ute = -1.613478125 lute = 9.48112101562515e-8
+ ua1 = 5.534185e-10 lua1 = -7.22371125000165e-19
+ ub1 = -4.333641125e-18 lub1 = 5.26789142906249e-25
+ uc1 = -2.8159131e-10 luc1 = 1.222685366175e-16 puc1 = -7.52316384526264e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.23 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.0e-05 wmax = 1.5e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.722382007957201+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.26470705697796e-07 wvth0 = -2.18005524689325e-06 pvth0 = 1.11019313448039e-12
+ k1 = 0.451376000000002 lk1 = 6.00222420000003e-8
+ k2 = 0.0527618062081521 lk2 = -6.41339581150145e-09 wk2 = -6.74947276007656e-08 pk2 = 3.43716900306898e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 50706.2890271588 lvsat = 0.00379987631291939 wvsat = -0.210762068777969 pvsat = 1.07330583525181e-7
+ ua = 1.18868819284835e-08 lua = -3.98065566078024e-15 wua = 4.71010489285566e-17 pua = -2.39862091668607e-23
+ ub = -9.66438145427305e-18 lub = 4.29465601563855e-24 wub = 1.47999308492692e-23 pub = -7.53686478499033e-30
+ uc = -1.43920874999999e-12 luc = -1.5724576940625e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0359168962159787 lu0 = -5.96917194798718e-09 wu0 = 5.57931960221544e-08 pu0 = -2.8412685074282e-14
+ a0 = 0.177126450000001 la0 = 3.202436703375e-7
+ keta = -0.1420657375 lketa = 2.2998105571875e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.123592234725+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 9.02619893870626e-9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.96298695527804+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.76447331197534e-06 wnfactor = -4.59795604474487e-05 pnfactor = 2.34150911578633e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.04625e-05 lcit = -1.0420528125e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.200224106952453 leta0 = 1.14038953215537e-07 weta0 = 5.87277493961004e-07 peta0 = -2.99071063799642e-13
+ etab = -0.0125364840599803 letab = 6.38420450754495e-09 wetab = 4.23712825280672e-07 petab = -2.15775756274182e-13
+ dsub = 0.42597171955 ldsub = -5.98739787258375e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.109122578548096 lpclm = 5.8962794299938e-07 wpclm = 1.30709898197858e-05 ppclm = -6.65640156572595e-12
+ pdiblc1 = 1.6849454761 lpdiblc1 = -5.69232019448926e-7
+ pdiblc2 = 0.00785230350750001 lpdiblc2 = -1.24879400639438e-9
+ pdiblcb = -0.025
+ drout = 0.857525935449999 ldrout = 1.72206730045879e-8
+ pscbe1 = 488447117.0 lpscbe1 = -51.4865790022495
+ pscbe2 = 1.539618939e-08 lpscbe2 = -3.72196255357505e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.19739062200001e-05 lalpha0 = 5.28379631080351e-11
+ alpha1 = 0.0
+ beta0 = 44.8934311524999 lbeta0 = 4.00699942758933e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.57161248473042e-08 lagidl = 1.10043398859897e-14 wagidl = 2.56064236488265e-13 pagidl = -1.30400712431649e-19
+ bgidl = 1557438821.0727 lbgidl = 76.2658803687245 wbgidl = 7617.61146653563 pbgidl = -0.00387926863933326
+ cgidl = -550.9458131622 lcgidl = 0.00039769665535285 wcgidl = 0.00638265358833322 pcgidl = -3.25036633985869e-9
+ egidl = 1.1826331595 legidl = -2.11731376402875e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.517158384853391 lkt1 = -1.22844417634105e-08 wkt1 = -8.0834718146496e-06 pkt1 = 4.11650802161031e-12
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.65197825000001 lute = 1.144173988125e-7
+ ua1 = 5.52e-10
+ ub1 = -7.96137600000001e-18 lub1 = 2.374213128e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.24 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.916781+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.0252804
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.704411452e-9
+ ub = -1.7524e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209856
+ a0 = 0.8967395
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1342734
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.1682+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.06764e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.622251
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.25 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.916781+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.59521
+ k2 = 0.0252804
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.704411452e-9
+ ub = -1.7524e-19
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0209856
+ a0 = 0.8967395
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1342734
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.1682+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.06764e-9
+ bgidl = 1704700000.0
+ cgidl = 700.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.622251
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.26 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.9182127628125+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.13241700247643e-8
+ k1 = 0.604152409375 lk1 = -7.07277513492169e-8
+ k2 = 0.02329948529375 lk2 = 1.56675496404078e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 297721.476875 lvsat = -0.772903590973594
+ ua = 2.44976570406838e-09 lua = 2.0140568818282e-15
+ ub = 8.85170975000002e-20 lub = -2.08612082340188e-24
+ uc = -5.15756313125e-11 luc = 9.17760209583907e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0202516383125 lu0 = 5.80508647685937e-9
+ a0 = 0.916541610412501 la0 = -1.56619841780065e-7
+ keta = -0.00495672689374999 lketa = -2.34839323906078e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1097586887125 lags = 1.9389298025066e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.094776478466875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.2431928936881e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.349198275+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.43156060654374e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.64831926658375 lpclm = 5.78838869829002e-06 ppclm = 3.23117426778526e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00455412315405625 lpdiblc2 = -1.27602734399944e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 562123300.169375 lpscbe1 = -1806.55551118713 ppscbe1 = 6.93889390390723e-18
+ pscbe2 = -1.5317388699625e-08 lpscbe2 = 2.39795383634009e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.815322348125e-05 lalpha0 = -2.17393918220826e-10
+ alpha1 = 0.0
+ beta0 = 39.1402881918125 lbeta0 = -6.91460005559311e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.57060410499999e-09 lagidl = -3.97806884747124e-15
+ bgidl = 1478354425.0 lbgidl = 1790.22373906875
+ cgidl = 932.600375000001 lcgidl = -0.00183969451596875
+ egidl = 1.20931880529938 legidl = -4.07967463450158e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.6304477199375 lkt1 = 6.4829907165672e-8
+ kt2 = -0.019032
+ at = 673047.845625 lat = -1.92232617300953
+ ute = -1.22055006875 lute = -1.31174856873906e-6
+ ua1 = 1.375495223e-09 lua1 = -5.29077591251275e-15
+ ub1 = -2.6104100625e-18 lub1 = -4.22820546317189e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.27 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.874172617125001+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.60839769504095e-7
+ k1 = 0.602594105000001 lk1 = -6.46359499712487e-8
+ k2 = 0.026832087675 lk2 = 1.8577237815062e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 84545.0750000001 lvsat = 0.06045625805625
+ ua = 3.31386607100375e-09 lua = -1.36392747761391e-15
+ ub = -1.45999138375e-18 lub = 3.96738595692469e-24 wub = -2.93873587705572e-39
+ uc = -5.4923007875e-11 luc = 1.04861752785344e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.020938342575 lu0 = 3.12058783868126e-9
+ a0 = 0.8237225450125 la0 = 2.06233089634885e-7
+ keta = -0.0050873285 lketa = -2.2973378061375e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.121306802125 lags = 1.48748517892844e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.064087020519875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.07540834542429e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.4583077875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.85809696828438e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0190949250000001 leta0 = 2.3809316444375e-7
+ etab = -0.1224012755 letab = 2.04849686248375e-7
+ dsub = 0.81474168125 ldsub = -9.95848917426563e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04876570365625 lpclm = -8.45940721620696e-7
+ pdiblc1 = 0.581562116725 lpdiblc1 = -7.48864204807207e-7
+ pdiblc2 = -0.001133342292 lpdiblc2 = 9.47345085500101e-9
+ pdiblcb = 0.165925 lpdiblcb = -7.4637355625e-07 wpdiblcb = -4.2351647362715e-22 ppdiblcb = -1.21169035041947e-27
+ drout = 0.139965000000001 ldrout = 1.64202182375e-6
+ pscbe1 = -156170353.9325 lpscbe1 = 1001.43395611063 ppscbe1 = -1.73472347597681e-18
+ pscbe2 = 7.6074691134375e-08 lpscbe2 = -1.17479104457055e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.4063189874125e-05 lalpha0 = -8.41274543421732e-11
+ alpha1 = -9.54625e-11 lalpha1 = 3.73186778125e-16
+ beta0 = 70.183410779125 lbeta0 = -0.000128269927030044
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.70826975625e-09 lagidl = -6.06988294620296e-16
+ bgidl = 2620002425 lbgidl = -2672.76370493125
+ cgidl = 455.747206250001 lcgidl = 2.44437339671881e-5
+ egidl = -1.5853225474425 legidl = 6.84527707370459e-06 wegidl = 1.6940658945086e-21 pegidl = 6.46234853557053e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.699418447125 lkt1 = 3.34453722423406e-7
+ kt2 = -0.019032
+ at = 210435.60875 lat = -0.113859286005937
+ ute = -1.7051169625 lute = 5.82544560653127e-7
+ ua1 = -4.84145456e-10 lua1 = 1.979024411868e-15 wua1 = -7.88860905221012e-31 pua1 = -1.88079096131566e-36
+ ub1 = -3.7199705125e-18 lub1 = 1.09343725990624e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.28 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.001397066+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 8.20635095105001e-8
+ k1 = 0.5590564875 lk1 = 1.84882462406245e-8
+ k2 = 0.023068907675 lk2 = 9.04257519650625e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 178330.86925 lvsat = -0.118604269615562
+ ua = 3.4633305675583e-09 lua = -1.64929256766068e-15
+ ub = 5.520602825e-19 lub = 1.25876313136875e-25
+ uc = 5.32329505e-13 luc = -1.01635010742125e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02660714225 lu0 = -7.70256794081251e-9
+ a0 = 1.02912416645 la0 = -1.85929956094663e-7
+ keta = 0.0443016559999999 lketa = -1.17269296718e-7
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.27952192815 lags = 9.14030771170387e-07 pags = -1.61558713389263e-27
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.15919953277725+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 7.40527294849646e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.574624755+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.70925138483748e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.454625e-05 lcit = -8.6799278125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.27451185329925 leta0 = -2.49561605911593e-7
+ etab = -0.028844949 letab = 2.622726987825e-8
+ dsub = 0.0649191575000003 ldsub = 4.35749736043125e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0624851574600003 lpclm = 1.0371154112045e-6
+ pdiblc1 = -0.00178611264999984 lpdiblc1 = 3.64893402127012e-7
+ pdiblc2 = 0.005940118645525 lpdiblc2 = -4.03155443996861e-9
+ pdiblcb = -0.40685 lpdiblcb = 3.471971125e-7
+ drout = 1.5358306539575 ldrout = -1.02303467606836e-6
+ pscbe1 = 430963245.09 lpscbe1 = -119.550867823082
+ pscbe2 = 1.4532757728e-08 lpscbe2 = 1.98318990660059e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.165892571425e-05 lalpha0 = 1.17722494844932e-10 walpha0 = -3.67127976680807e-26 palpha0 = -1.66222800528309e-31
+ alpha1 = 1.90925e-10 lalpha1 = -1.7359855625e-16
+ beta0 = -39.87379705625 lbeta0 = 8.18567970296454e-05 wbeta0 = -5.42101086242752e-20 pbeta0 = -1.03397576569128e-25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.0118678375e-09 lagidl = -1.18663293124687e-15
+ bgidl = 793843600.000001 lbgidl = 813.8300317
+ cgidl = 559.9750875 lcgidl = -0.000174553348309375
+ egidl = 3.11021319877 legidl = -2.11967454975162e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.73964705275 lkt1 = 4.11260187712937e-7
+ kt2 = -0.019032
+ at = 260637.4 lat = -0.20970705595
+ ute = -1.3447176 lute = -1.05547922200001e-7
+ ua1 = 5.524e-10
+ ub1 = -3.72798415e-18 lub1 = 1.24643763387503e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.29 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.876262085+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -3.1715471963749e-8
+ k1 = 0.590241525000001 lk1 = -9.86674910624936e-9
+ k2 = 0.02128655125 lk2 = 1.06631827759375e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8367.10762500018 lvsat = 0.0359352806419687
+ ua = -8.27123482416499e-10 lua = 2.2518027772789e-15
+ ub = 3.741906275e-18 lub = -2.77449115554375e-24
+ uc = 6.082695725e-12 luc = -6.06302059295625e-18 wuc = -1.23259516440783e-32 puc = -5.87747175411144e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.01445975725 lu0 = 3.34244187043749e-9
+ a0 = 0.757708623749998 la0 = 6.08546261053134e-8
+ keta = -0.1537600425 lketa = 6.2818302643125e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.74210549 lags = -1.4883958782501e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.095254583405+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.59107842682463e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.855709525+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.33575146560625e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.273125e-05 lcit = 1.61221390625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.039032375e-05 leta0 = 4.77441026196875e-11
+ etab = 0.0007545356125 letab = -6.86061505665625e-10
+ dsub = 1.499306975 ldsub = -8.68467387018751e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.0219588243125 lpclm = -7.44536020381139e-7
+ pdiblc1 = 0.1958620354125 lpdiblc1 = 1.85181823501184e-7
+ pdiblc2 = -0.033618504135125 lpdiblc2 = 3.19371233233374e-08 wpdiblc2 = -5.29395592033938e-23 ppdiblc2 = 1.26217744835362e-29
+ pdiblcb = -0.025
+ drout = 0.335842470275 ldrout = 6.80545799449566e-8
+ pscbe1 = -56987686.124999 lpscbe1 = 324.118516384156
+ pscbe2 = 1.82815146225e-08 lpscbe2 = -3.38872530725814e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0002471576267875 lalpha0 = -1.63068955517284e-10
+ alpha1 = 0.0
+ beta0 = 67.1968940187498 lbeta0 = -1.54972288302984e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.50369049999999e-09 lagidl = 1.2011638487125e-14
+ bgidl = 1269024000 lbgidl = 381.772252999999
+ cgidl = -171.03 lcgidl = 0.000490113027499999
+ egidl = 1.8355566512875 legidl = -9.6069308395316e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.0223996624999998 lkt1 = -2.40897001871876e-7
+ kt2 = -0.019032
+ at = 47731.2499999999 lat = -0.0161221390625
+ ute = -1.39342125 lute = -6.12641284375002e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.30 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.794303062499997+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -8.98449086718744e-8
+ k1 = 0.5943829125 lk1 = -1.28040281906251e-8
+ k2 = 0.0265255762499999 lk2 = 6.94740429468747e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 61237.988625 lvsat = -0.00156339170728126
+ ua = -2.037867569625e-09 lua = 3.11052302113153e-15
+ ub = 2.53193054975e-18 lub = -1.91631587241019e-24 wub = 5.87747175411144e-39 pub = -1.40129846432482e-45
+ uc = 2.7825305e-12 luc = -3.722378407125e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00638258624999999 lu0 = 9.0711754021875e-9
+ a0 = 0.9390707625 la0 = -6.77764708031244e-8
+ keta = 0.0155643187500001 lketa = -5.72750005734375e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.625540699999998 lags = 9.55119101474999e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '0.01132308791625+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.96794291163503e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.1799136+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -8.56443205800002e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0601722599225 leta0 = 4.27175501155331e-08 weta0 = -5.21123785908407e-23 peta0 = -7.37584946381646e-29
+ etab = -0.0007545356125 letab = 3.84247260665625e-10
+ dsub = 0.189319827725 ldsub = 6.06409971860439e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.221698298187498 lpclm = 5.32298757773016e-7
+ pdiblc1 = 0.1763525393125 lpdiblc1 = 1.99018933610109e-7
+ pdiblc2 = 0.0267160385535 lpdiblc2 = -1.08551510785699e-8
+ pdiblcb = -0.025
+ drout = -0.738324518225 ldrout = 8.29907516538581e-7
+ pscbe1 = 432224423.35 lpscbe1 = -22.8551722609873
+ pscbe2 = 1.054562873625e-08 lpscbe2 = 2.09795175756469e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.00012163830041875 lalpha0 = 9.84995558537484e-11 walpha0 = -2.06795153138257e-25 palpha0 = 1.97215226305253e-31
+ alpha1 = 0.0
+ beta0 = 26.4659450524999 lbeta0 = 1.33911967240144e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.84437134625e-08 lagidl = -6.39155777327812e-15
+ bgidl = 2062179625.0 lbgidl = -180.773374031251
+ cgidl = 1258.4125 lcgidl = -0.000523719065625
+ egidl = -0.246745445500001 legidl = 5.16179678193375e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.0943169337500001 lkt1 = -3.23678247762187e-7
+ kt2 = -0.019032
+ at = 42823.75 lat = -0.0126414946875
+ ute = -1.613478125 lute = 9.48112101562515e-8
+ ua1 = 5.534185e-10 lua1 = -7.22371125000165e-19
+ ub1 = -4.333641125e-18 lub1 = 5.26789142906252e-25
+ uc1 = -2.8159131e-10 luc1 = 1.222685366175e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.31 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7e-06 wmax = 1.0e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.839765803011765+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -6.66930080662589e-08 wvth0 = -1.00909953805139e-06 pvth0 = 5.13883939752668e-13
+ k1 = 0.451376000000002 lk1 = 6.00222420000003e-8
+ k2 = 0.0469472870918334 lk2 = -3.4523519515161e-09 wk2 = -9.49230613996067e-09 pk2 = 4.83395690177486e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8589.48890543205 lvsat = 0.0252478567749088 wvsat = 0.209371796529108 pvsat = -1.06622587382449e-7
+ ua = 1.19027771371721e-08 lua = -3.98875029580488e-15 wua = -1.1146074700276e-16 pua = 5.67613854111454e-23
+ ub = -8.63997172801878e-18 lub = 3.77297536254356e-24 wub = 4.58098694314493e-24 pub = -2.33286760079656e-30
+ uc = -1.43920874999999e-12 luc = -1.5724576940625e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0377341307796053 lu0 = -6.89459864951403e-09 wu0 = 3.7665470763363e-08 pu0 = -1.91811409862427e-14
+ a0 = 0.177126449999999 la0 = 3.202436703375e-7
+ keta = -0.1420657375 lketa = 2.29981055718751e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.123592234725+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 9.02619893870626e-9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.28643936341503+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 1.07808549180894e-07 wnfactor = -9.30435847838924e-06 pnfactor = 4.73824455511974e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.04625e-05 lcit = -1.0420528125e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.011003604573435 leta0 = 6.47124112097818e-09 weta0 = -1.51981313606907e-06 peta0 = 7.73964839543175e-13
+ etab = 0.0629137474333006 letab = -3.20388258804083e-08 wetab = -3.2893688466805e-07 petab = 1.67511108517205e-13
+ dsub = 0.425971719550001 ldsub = -5.98739787258381e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.43696958545631 lpclm = -5.95828145268627e-07 wpclm = -1.01503222938887e-05 ppclm = 5.16905162816281e-12
+ pdiblc1 = 1.6849454761 lpdiblc1 = -5.69232019448926e-7
+ pdiblc2 = 0.00785230350750001 lpdiblc2 = -1.24879400639437e-9
+ pdiblcb = -0.025
+ drout = 0.857525935449999 ldrout = 1.72206730045871e-8
+ pscbe1 = 488447117.0 lpscbe1 = -51.4865790022504
+ pscbe2 = 1.539618939e-08 lpscbe2 = -3.72196255357505e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.19739062200001e-05 lalpha0 = 5.28379631080351e-11
+ alpha1 = 0.0
+ beta0 = 44.8934311524999 lbeta0 = 4.00699942758933e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.60424053956415e-08 lagidl = -5.16869164023044e-15 wagidl = -6.0741266989607e-14 pagidl = 3.09324902144574e-20
+ bgidl = 2321075000.0 lbgidl = -312.61584375
+ cgidl = -772.087304690801 lcgidl = 0.000510312959913791 wcgidl = 0.00858863859543624 pcgidl = -4.37376420472591e-9
+ egidl = 1.1826331595 legidl = -2.11731376402875e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 1.01040992042532 lkt1 = -7.90198601226594e-07 wkt1 = -2.33216469552689e-05 pkt1 = 1.18765487119707e-11
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.65197825 lute = 1.144173988125e-7
+ ua1 = 5.52e-10
+ ub1 = -7.961376e-18 lub1 = 2.374213128e-24
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.32 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.905854920584+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = -7.62142769580179e-8
+ k1 = 0.59521
+ k2 = 0.0256978399194 wk2 = -2.91182961601904e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70511538307553e-09 wua = -4.91023320506719e-18
+ ub = -3.724600519e-20 wub = -9.62569659121435e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0221657757912 wu0 = -8.23225250202285e-9
+ a0 = 0.896182001275701 wa0 = 3.88880224642466e-9
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1361319778533 wags = -1.29644094524902e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.8729719259+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = -4.91609851143144e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.04819616582e-09 wagidl = 4.19883054153556e-14
+ bgidl = 1704700000.0
+ cgidl = -46.3169000000003 wcgidl = 0.0052058932348374
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.0645073236570002 wkt1 = -4.79044560171993e-6
+ kt2 = -0.019032
+ at = 383230.8076 wat = 0.32623597604981
+ ute = -1.0139878669 wute = -2.59774072418386e-6
+ ua1 = 2.409316835472e-09 wua1 = -1.18774883569658e-14
+ ub1 = -1.8571058029e-18 wub1 = -8.9836364255844e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.33 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.905854920584+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = -7.62142769580179e-8
+ k1 = 0.59521
+ k2 = 0.0256978399194 wk2 = -2.91182961601915e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.70511538307553e-09 wua = -4.91023320506719e-18
+ ub = -3.72460051900002e-20 wub = -9.62569659121435e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0221657757912 wu0 = -8.23225250202285e-9
+ a0 = 0.8961820012757 wa0 = 3.88880224642466e-9
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1361319778533 wags = -1.29644094524906e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.8729719259+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = -4.91609851143144e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.04819616582001e-09 wagidl = 4.19883054153555e-14
+ bgidl = 1704700000.0
+ cgidl = -46.3168999999989 wcgidl = 0.0052058932348374
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.0645073236570002 wkt1 = -4.79044560171992e-6
+ kt2 = -0.019032
+ at = 383230.8076 wat = 0.326235976049809
+ ute = -1.0139878669 wute = -2.59774072418387e-6
+ ua1 = 2.409316835472e-09 wua1 = -1.18774883569658e-14
+ ub1 = -1.8571058029e-18 wub1 = -8.9836364255844e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.34 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.939506042855864+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 2.66155138828752e-07 wvth0 = 1.48530125105373e-07 pvth0 = -1.7775596620199e-12
+ k1 = 0.604152409375 lk1 = -7.07277513492185e-8
+ k2 = 0.0233233005303496 lk2 = 1.87808256628471e-08 wk2 = -1.66121896877705e-10 pk2 = -2.17164887776193e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 358260.418207494 lvsat = -1.25172121270762 wvsat = -0.422286116161978 pvsat = 3.33996646425413e-6
+ ua = 2.45066693860442e-09 lua = 2.01249635943307e-15 wua = -6.28651283955156e-18 pua = 1.08853396991537e-23
+ ub = 2.20141131414774e-19 lub = -2.03573921019131e-24 wub = -9.18136340874673e-25 pub = -3.51434222343205e-31
+ uc = -5.15756313125e-11 luc = 9.17760209583907e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0214357041561551 lu0 = 5.77431907947882e-09 wu0 = -8.25938735286063e-09 pu0 = 2.14616318988171e-16
+ a0 = 0.919712726966413 la0 = -1.86110392169274e-07 wa0 = -2.21199522815272e-08 pa0 = 2.05709741750216e-13
+ keta = -0.00495672689375 lketa = -2.34839323906078e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0938470206943461 lags = 3.34442297409455e-07 wags = 1.10990981030558e-07 pags = -9.80394172178052e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.094776478466875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.24319289368818e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.31704838893699+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 4.39693823472468e-06 wnfactor = 2.24259794138652e-07 pnfactor = -4.06563789283305e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.64831926658375 lpclm = 5.78838869829003e-06 wpclm = -4.2351647362715e-22 ppclm = -4.8467614016779e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00455412315405625 lpdiblc2 = -1.27602734399944e-08 wpdiblc2 = 1.32348898008484e-23
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 562123300.169375 lpscbe1 = -1806.55551118713
+ pscbe2 = -1.5317388699625e-08 lpscbe2 = 2.39795383634009e-13 ppscbe2 = 3.85185988877447e-34
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.815322348125e-05 lalpha0 = -2.17393918220827e-10
+ alpha1 = 0.0
+ beta0 = 39.1402881918125 lbeta0 = -6.9146000555929e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.21755219505243e-08 lagidl = 1.04589692511696e-13 wagidl = 1.37738036009503e-13 pagidl = -7.5730855670176e-19
+ bgidl = 1297223857.55941 lbgidl = 3222.83067959827 wbgidl = 1263.46649213122 pbgidl = -0.00999307235288885
+ cgidl = -61.7073690126253 lcgidl = 0.000121727067038106 wcgidl = 0.00693573997574189 pcgidl = -1.36817903354989e-8
+ egidl = 1.20931880529937 legidl = -4.07967463450159e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.192931677225396 lkt1 = -1.01574031846084e-06 wkt1 = -5.74343852242234e-06 pkt1 = 7.53745925806556e-12
+ kt2 = -0.019032
+ at = 712808.007523131 lat = -2.60670846849202 wat = -0.277344862271669 pat = 4.77387174549415e-6
+ ute = -0.484174902819705 lute = -4.19042318615206e-06 wute = -5.1365452056878e-06 pute = 2.00800393453351e-11
+ ua1 = 4.74237759823923e-09 lua1 = -1.84527608379167e-14 wua1 = -2.3485506196833e-14 pua1 = 9.18107150999694e-20
+ ub1 = -5.12655569903866e-19 lub1 = -1.06335930053247e-23 wub1 = -1.46327731843617e-23 pub1 = 4.46804349093595e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.35 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.825665150885932+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.78877368104704e-07 wvth0 = -3.38361211347436e-07 pvth0 = 1.2582029500826e-13
+ k1 = 0.602594105 lk1 = -6.46359499712495e-8
+ k2 = 0.0274254924827725 lk2 = 2.74433177283797e-09 wk2 = -4.13926319275697e-09 pk2 = -6.18448616670344e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -12784.3819762375 lvsat = 0.198785672410632 wvsat = 0.678916371347068 pvsat = -9.64909360040613e-7
+ ua = 3.30616298981007e-09 lua = -1.33185157874259e-15 wua = 5.37324269001763e-17 pua = -2.23743700478361e-22
+ ub = -1.19286643284898e-18 lub = 3.48806061040679e-24 wub = -1.86331567026269e-24 pub = 3.34350807106689e-30
+ uc = -5.4923007875e-11 luc = 1.04861752785344e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0223473675748525 lu0 = 2.2103988599361e-09 wu0 = -9.82857779912106e-09 pu0 = 6.34897407103223e-15
+ a0 = 0.801686911444114 la0 = 2.7528202716127e-07 wa0 = 1.53708372032056e-07 pa0 = -4.81647135072676e-13
+ keta = -0.0050873285 lketa = -2.2973378061375e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.146165515536263 lags = 1.29916221448692e-07 wags = -1.7340061302974e-07 pags = 1.31363666902172e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0640870205198749+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.07540834542429e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '6.4053761868607+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -3.76685720930859e-06 wnfactor = -1.3581670478047e-05 pnfactor = 1.33144539882114e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0190949249999999 leta0 = 2.3809316444375e-7
+ etab = -0.1224012755 letab = 2.04849686248375e-7
+ dsub = 0.81474168125 ldsub = -9.95848917426562e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04876570365625 lpclm = -8.45940721620694e-07 wpclm = -3.3881317890172e-21
+ pdiblc1 = 0.581562116725 lpdiblc1 = -7.48864204807207e-7
+ pdiblc2 = -0.001133342292 lpdiblc2 = 9.47345085500101e-09 ppdiblc2 = -1.26217744835362e-29
+ pdiblcb = 0.165925 lpdiblcb = -7.4637355625e-07 wpdiblcb = 2.11758236813575e-22 ppdiblcb = 2.01948391736579e-28
+ drout = 0.139965 ldrout = 1.64202182375e-6
+ pscbe1 = -156170353.9325 lpscbe1 = 1001.43395611063 ppscbe1 = 8.67361737988404e-19
+ pscbe2 = 7.6074691134375e-08 lpscbe2 = -1.17479104457056e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.4063189874125e-05 lalpha0 = -8.41274543421732e-11
+ alpha1 = -9.54625e-11 lalpha1 = 3.73186778125e-16
+ beta0 = 70.183410779125 lbeta0 = -0.000128269927030044
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.3145748246658e-08 lagidl = 5.60251699336144e-15 wagidl = -4.49042835860022e-14 pagidl = -4.33140688230312e-20
+ bgidl = 2982263559.88119 lbgidl = -3364.41077670316 wbgidl = -2526.93298426244 pbgidl = 0.00482454680020307
+ cgidl = -507.04077638725 lcgidl = 0.00186264668981736 wcgidl = 0.00671587558233508 pcgidl = -1.28222854555732e-8
+ egidl = -1.5853225474425 legidl = 6.84527707370459e-06 pegidl = -9.69352280335579e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.209402020212483 lkt1 = -1.08012700678311e-06 wkt1 = -6.33942809360739e-06 pkt1 = 9.86733148922069e-12
+ kt2 = -0.019032
+ at = -163282.090709361 lat = 0.818146748023348 wat = 2.606847631823 pat = -6.50115776204545e-6
+ ute = -1.82338412242998 lute = 1.04488045560938e-06 wute = 8.24966187664906e-07 pute = -3.22499906912903e-12
+ ua1 = -4.84145456e-10 lua1 = 1.979024411868e-15 wua1 = 4.93038065763132e-31 pua1 = 2.63310734584192e-36
+ ub1 = -2.65182721204045e-18 lub1 = -2.27103626330222e-24 wub1 = -7.45077591261736e-24 pub1 = 1.66042120747928e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.36 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.98308130697379+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.21669427906037e-07 wvth0 = -1.27760588036333e-07 pvth0 = -2.76268945048482e-13
+ k1 = 0.5590564875 lk1 = 1.8488246240625e-8
+ k2 = 0.0202297791236843 lk2 = 1.64827475036771e-08 wk2 = 1.98041878967608e-08 pk2 = -5.18985201593654e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 130834.0178725 lvsat = -0.0754177575005706 wvsat = 0.331311721953777 pvsat = -3.01245183186472e-7
+ ua = 3.48199372939773e-09 lua = -1.66755641830033e-15 wua = -1.30183877600178e-16 pua = 1.27398503888937e-22
+ ub = 1.41860159332835e-18 lub = -1.49788471857228e-24 wub = -6.04451212045235e-24 pub = 1.13264573935915e-29
+ uc = 5.32329505000001e-13 luc = -1.01635010742125e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0298784458896418 lu0 = -1.21683124125754e-08 wu0 = -2.28188018879247e-08 pu0 = 3.11505594125803e-14
+ a0 = 1.06570133789856 la0 = -2.28787516546874e-07 wa0 = -2.5514208427216e-07 pa0 = 2.98950598626143e-13
+ keta = 0.0443016560000001 lketa = -1.17269296718e-07 pketa = 2.01948391736579e-28
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.235271615490397 lags = 8.58175063861341e-07 wags = -3.0866566644018e-07 pags = 3.89618470126057e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.196533217860814+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.45332067730759e-07 wvoff = 2.60419104281404e-07 pvoff = -4.97205174849272e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.62704043431987+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -3.7156967377e-07 wnfactor = -7.34106874064903e-06 pnfactor = 1.39958512108437e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.454625e-05 lcit = -8.6799278125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.275607482161874 leta0 = -2.51653435317558e-07 weta0 = -7.64249996727589e-09 peta0 = 1.45914430625213e-14
+ etab = -0.028844949 letab = 2.622726987825e-8
+ dsub = -0.489646099812167 ldsub = 1.49455345356638e-06 wdsub = 3.86834000585713e-06 pdsub = -7.38562815618273e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0624851574599994 lpclm = 1.03711541120449e-6
+ pdiblc1 = -0.00178611265000006 lpdiblc1 = 3.64893402127012e-7
+ pdiblc2 = 0.005940118645525 lpdiblc2 = -4.0315544399686e-9
+ pdiblcb = -0.40685 lpdiblcb = 3.471971125e-7
+ drout = 1.5358306539575 ldrout = -1.02303467606836e-6
+ pscbe1 = 430963245.09 lpscbe1 = -119.550867823082
+ pscbe2 = 1.4532757728e-08 lpscbe2 = 1.98318990660059e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.165892571425e-05 lalpha0 = 1.17722494844932e-10 walpha0 = -9.01944115984444e-26 palpha0 = -1.40465744471283e-31
+ alpha1 = 1.90925e-10 lalpha1 = -1.7359855625e-16
+ beta0 = -39.87379705625 lbeta0 = 8.18567970296453e-05 pbeta0 = 7.75481824268463e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.83690786984924e-08 lagidl = -4.37012667180351e-15 wagidl = -7.92216110714661e-14 pagidl = 2.22062886785908e-20
+ bgidl = 510872136.567474 lbgidl = 1354.09329825855 wbgidl = 1973.85216271455 pbgidl = -0.00376857724166276
+ cgidl = 559.9750875 lcgidl = -0.000174553348309375
+ egidl = 3.11021319877 legidl = -2.11967454975162e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.14541453851815 lkt1 = 1.50655650797336e-06 wkt1 = 2.83040918553153e-06 pkt1 = -7.6401803359753e-12
+ kt2 = -0.019032
+ at = 479122.9163365 lat = -0.408365011678963 wat = -1.52403392098737 pat = 1.38572784265777e-6
+ ute = -1.10818328014005 lute = -3.2061675253266e-07 wute = -1.64993237532981e-06 pute = 1.50020101226863e-12
+ ua1 = 5.524e-10
+ ub1 = -4.06901154289045e-18 lub1 = 4.34722920373141e-25 wub1 = 2.37881816362812e-24 pub1 = -2.16294041527887e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.37 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.450441033032307+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -3.62633741175256e-07 wvth0 = -2.97029175366384e-06 pvth0 = 2.30830251729832e-12
+ k1 = 0.590241525 lk1 = -9.86674910625021e-9
+ k2 = 0.0424658276553063 lk2 = -3.73537962370024e-09 wk2 = -1.47734898884288e-07 pk2 = 1.00436394496303e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6473.00539822539 lvsat = 0.0376574930916637 wvsat = 0.0132122078013457 pvsat = -1.20131999433738e-8
+ ua = -7.9321575854206e-10 lua = 2.21967780860892e-15 wua = -2.36521496869073e-16 pua = 2.2408598420913e-22
+ ub = -8.00767241092021e-19 lub = 5.20076394124436e-25 wub = 3.168717380713e-23 pub = -2.29810780360628e-29
+ uc = 6.082695725e-12 luc = -6.06302059295625e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00396046101905728 lu0 = 1.13976153310036e-08 wu0 = 7.32372738969444e-08 pu0 = -5.6188427494812e-14
+ a0 = 0.709709787186945 la0 = 9.48978009376614e-08 wa0 = 3.34813292508427e-07 pa0 = -2.37466327711596e-13
+ keta = -0.1537600425 lketa = 6.28183026431251e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.663999937383494 lags = 4.0512404410758e-08 wags = 5.44821064576605e-07 pags = -3.8641434005096e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '0.091413842012819+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.16483796459342e-07 wvoff = -1.30209552140702e-06 pvoff = 9.2351124855793e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '10.5414557000471+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.74925175413252e-06 wnfactor = -3.96606154137479e-05 pnfactor = 3.07861329335995e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.273125e-05 lcit = 1.61221390625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.000286792136043527 leta0 = -1.31809791157168e-09 weta0 = -2.07298020043692e-09 peta0 = 9.52735721452314e-15
+ etab = -0.00206103367336456 letab = 1.87399486750673e-09 wetab = 1.96398515128068e-08 petab = -1.78575349880196e-14
+ dsub = 4.27216422708862 ldsub = -2.83512258616816e-06 wdsub = -1.93419160276526e-05 pdsub = 1.3718297142286e-11
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.0219588243125 lpclm = -7.4453602038114e-7
+ pdiblc1 = 0.1958620354125 lpdiblc1 = 1.85181823501185e-7
+ pdiblc2 = -0.033618504135125 lpdiblc2 = 3.19371233233374e-08 ppdiblc2 = -3.78653234506086e-29
+ pdiblcb = -0.025
+ drout = 0.335842470275001 ldrout = 6.80545799449558e-8
+ pscbe1 = -56987686.125 lpscbe1 = 324.118516384156
+ pscbe2 = 1.82815146225e-08 lpscbe2 = -3.38872530725811e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0002471576267875 lalpha0 = -1.63068955517284e-10 walpha0 = 8.27180612553028e-25
+ alpha1 = 0.0
+ beta0 = 67.19689401875 lbeta0 = -1.54972288302984e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.09421604184736e-08 lagidl = -6.70970122569643e-15 wagidl = -1.98422497005863e-13 pagidl = 1.30589694214441e-19
+ bgidl = 2683881317.16262 lbgidl = -621.715299197593 wbgidl = -9869.26081357275 pbgidl = 0.00699977323202648
+ cgidl = -171.03 lcgidl = 0.000490113027500001
+ egidl = 1.8355566512875 legidl = -9.60693083953159e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 5.14299323044094 lkt1 = -4.2111782559527e-06 wkt1 = -3.60309191934933e-05 pkt1 = 2.76944824926531e-11
+ kt2 = -0.019032
+ at = 47731.2500000001 lat = -0.0161221390625
+ ute = -1.39342125 lute = -6.12641284375002e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.38 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.938826503017104+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.62463465885398e-08 wvth0 = 1.00811545506126e-06 pvth0 = -5.13382795489948e-13
+ k1 = 0.5943829125 lk1 = -1.28040281906251e-8
+ k2 = 0.0296397732041287 lk2 = 5.36149949579745e-09 wk2 = -2.17229126868893e-08 pk2 = 1.10623932857985e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 63132.0908517746 lvsat = -0.0025279632662662 wvsat = -0.0132122078013461 pvsat = 6.72831682283543e-9
+ ua = -2.07824714718519e-09 lua = 3.13108632100405e-15 wua = 2.81665562773846e-16 pua = -1.43438187842588e-22
+ ub = 2.89531234164961e-18 lub = -2.10136804993507e-24 wub = -2.53475006677899e-24 pub = 1.2908214715072e-30
+ uc = 2.7825305e-12 luc = -3.722378407125e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00942532429384987 lu0 = 7.52166105335693e-09 wu0 = -2.12244549170204e-08 pu0 = 1.08085536664926e-14
+ a0 = 0.9390707625 la0 = -6.77764708031261e-8
+ keta = 0.0155643187500001 lketa = -5.72750005734375e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.6255407 lags = 9.55119101475e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '0.01132308791625+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.96794291163503e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.27548953062954+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 1.1338475152691e-07 wnfactor = 1.32842072569939e-05 pnfactor = -6.76498254562417e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.065947586695414 leta0 = 4.56586352746396e-08 weta0 = 4.02854800368163e-08 peta0 = -2.05153807087487e-14
+ etab = 0.00206103367336456 letab = -1.0495813981609e-09 wetab = -1.96398515128068e-08 petab = 1.00015943828969e-14
+ dsub = 0.189288862197213 ldsub = 6.06567663810691e-08 wdsub = 2.15998366941687e-10 pdsub = -1.09997168365768e-16
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2216982981875 lpclm = 5.32298757773016e-7
+ pdiblc1 = 0.1763525393125 lpdiblc1 = 1.99018933610109e-7
+ pdiblc2 = 0.0267160385535 lpdiblc2 = -1.08551510785699e-8
+ pdiblcb = -0.025
+ drout = -0.738324518224999 ldrout = 8.29907516538581e-7
+ pscbe1 = 432224423.35 lpscbe1 = -22.8551722609873
+ pscbe2 = 1.054562873625e-08 lpscbe2 = 2.09795175756471e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.00012163830041875 lalpha0 = 9.84995558537484e-11 palpha0 = 9.86076131526265e-32
+ alpha1 = 0.0
+ beta0 = 26.4659450525 lbeta0 = 1.33911967240144e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.571311371803e-08 lagidl = -1.00934998534068e-14 wagidl = -5.07073089348358e-14 pagidl = 2.58226970750651e-20
+ bgidl = 2062179625 lbgidl = -180.773374031251
+ cgidl = 1258.4125 lcgidl = -0.000523719065625
+ egidl = -0.2467454455 legidl = 5.16179678193375e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.4393147900623 lkt1 = 4.57323707589227e-07 wkt1 = 1.06977652733396e-05 pkt1 = -5.4478369654482e-12
+ kt2 = -0.019032
+ at = 42823.75 lat = -0.0126414946875
+ ute = -1.613478125 lute = 9.48112101562498e-8
+ ua1 = 5.534185e-10 lua1 = -7.22371125000165e-19
+ ub1 = -4.333641125e-18 lub1 = 5.26789142906249e-25
+ uc1 = -2.8159131e-10 luc1 = 1.222685366175e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.39 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.37663231406486+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 2.06706262687528e-07 wvth0 = 2.73578381900786e-06 pvth0 = -1.39319790982975e-12
+ k1 = 0.332563655574575 lk1 = 1.20527428398648e-07 wk1 = 8.28769092672963e-07 pk1 = -4.22050660443704e-13
+ k2 = 0.0418805836785902 lk2 = -8.72133238321973e-10 wk2 = 2.5850209917134e-08 pk2 = -1.31642194003004e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 102283.153988712 lvsat = -0.0224656421687514 wvsat = -0.444183304801394 pvsat = 2.2620034797011e-7
+ ua = 1.87124330232666e-08 lua = -7.4565675557985e-15 wua = -4.7611847659037e-14 pua = 2.42463334203646e-20
+ ub = -8.79517665810563e-18 lub = 3.85201347319029e-24 wub = 5.66361055189958e-24 pub = -2.88419367355486e-30
+ uc = -4.79277200709405e-11 luc = 2.21018166961265e-17 wuc = 3.24278100339609e-16 puc = -1.65138622597946e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0688744914242333 lu0 = -2.27528273077908e-08 wu0 = -1.79552433333764e-07 pu0 = 9.14370766752194e-14
+ a0 = -1.46008118556577 la0 = 1.15399165874937e-06 wa0 = 1.14202534526767e-05 pa0 = -5.81576407077563e-12
+ keta = -0.037954766283685 lketa = -3.00204065200334e-08 wketa = -7.2622045772696e-07 pketa = 3.69827768097455e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.44347029220031+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.71924099708008e-07 wvoff = 2.23129211650392e-06 pvoff = -1.13628551032962e-12
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '-5.69155831195651+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 4.17060386536385e-06 wnfactor = 4.63457334942904e-05 pnfactor = -2.36015647819674e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.04625e-05 lcit = -1.0420528125e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.61134784136532 leta0 = 3.23403714965289e-07 weta0 = 2.82136576809864e-06 peta0 = -1.43678051740423e-12
+ etab = -0.0491842326301592 letab = 2.50470704669086e-08 wetab = 4.5299652197369e-07 petab = -2.30688478815102e-13
+ dsub = 0.536120536598492 ldsub = -1.15967263807782e-07 wdsub = -7.68337125285635e-07 pdsub = 3.91275681051709e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.570174338286741 lpclm = 9.35559897897524e-07 wpclm = 1.08258477604091e-05 ppclm = -5.51306297198834e-12
+ pdiblc1 = 2.68942229835588 lpdiblc1 = -1.08076184118273e-06 wpdiblc1 = -7.00667383189752e-06 ppdiblc1 = 3.56814864889381e-12
+ pdiblc2 = 0.0401093439324827 lpdiblc2 = -1.76756918428168e-08 wpdiblc2 = -2.25007243604284e-07 ppdiblc2 = 1.14584938805482e-13
+ pdiblcb = -0.025
+ drout = -0.943896140671598 ldrout = 9.34594865269511e-07 wdrout = 1.25657224151941e-05 pdrout = -6.39909413993759e-12
+ pscbe1 = 29721003.5986633 lpscbe1 = 182.11969424738 wpscbe1 = 3199.8192328209 ppscbe1 = -0.00162950794431405
+ pscbe2 = 1.51162422576379e-08 lpscbe2 = -2.296331782021e-16 wpscbe2 = 1.95275610464662e-15 ppscbe2 = -9.94441046291318e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000572116254996407 lalpha0 = 3.2790545422242e-10 walpha0 = 3.76773378620299e-09 palpha0 = -1.91871843062387e-15
+ alpha1 = 0.0
+ beta0 = 2.63744925086473 lbeta0 = 2.55258582109971e-05 wbeta0 = 0.000294754319931834 pbeta0 = -1.50103637425286e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.54208791186093e-08 lagidl = -1.50371793836518e-14 wagidl = -1.95914764006587e-13 pagidl = 9.97695935703547e-20
+ bgidl = 3487818330.8615 lbgidl = -906.77988499122 wbgidl = -8138.55510028452 pbgidl = 0.00414455918481989
+ cgidl = 2760.087441315 lcgidl = -0.00128844702948966 wcgidl = -0.016049855607891 pcgidl = 8.17338896831847e-9
+ egidl = 1.27487022659837 legidl = -2.58703102822717e-07 wegidl = -6.43394680743017e-07 pegidl = 3.27648741168382e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -6.94299218526389 lkt1 = 3.26007142109564e-06 wkt1 = 3.21568799492525e-05 pkt1 = -1.63758911141568e-11
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.65197825 lute = 1.14417398812502e-7
+ ua1 = 5.52e-10
+ ub1 = -1.5434234681085e-17 lub1 = 6.17976641134254e-24 wub1 = 5.21265221955397e-23 pub1 = -2.65454314280786e-29
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.40 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.934970143102+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = 6.86469404582746e-8
+ k1 = 0.59521
+ k2 = 0.0253484040955 wk2 = -1.17323054373906e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.78879880790487e-09 wua = -4.21272594538509e-16
+ ub = -2.7812373201e-19 wub = 2.35904463274226e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0216317529636 wu0 = -5.57525076053175e-9
+ a0 = 0.5363746550628 wa0 = 1.79409082373201e-6
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0950869594429 wags = 1.91252863217461e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.2556405716+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = -1.84459969400494e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.52019415876e-08 wagidl = -2.84328906284581e-14
+ bgidl = 1599071667.0 wbgidl = 525.548066911517
+ cgidl = 1000.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.77537944851 wkt1 = -6.11634320688714e-7
+ kt2 = -0.019032
+ at = 448800.0
+ ute = -1.5361
+ ua1 = 2.2096e-11
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.41 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.934970143102+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = 6.86469404582746e-8
+ k1 = 0.59521
+ k2 = 0.0253484040955 wk2 = -1.17323054373911e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200000.0
+ ua = 2.78879880790487e-09 wua = -4.21272594538518e-16
+ ub = -2.7812373201e-19 wub = 2.35904463274226e-25
+ uc = -3.9972e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0216317529636 wu0 = -5.57525076053177e-9
+ a0 = 0.5363746550628 wa0 = 1.79409082373201e-6
+ keta = -0.0079259
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0950869594429 wags = 1.91252863217461e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.093204657+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.2556405716+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = -1.84459969400493e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.08353125
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 333712830.0
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.52019415876e-08 wagidl = -2.84328906284581e-14
+ bgidl = 1599071667.0 wbgidl = 525.548066911517
+ cgidl = 1000.0
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.77537944851 wkt1 = -6.11634320688714e-7
+ kt2 = -0.019032
+ at = 448800.0
+ ute = -1.5361
+ ua1 = 2.2096e-11
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.42 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.923219379389274+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -9.2939727894877e-08 wvth0 = 6.7496710507177e-08 pvth0 = 9.09745624071843e-15
+ k1 = 0.604152409375 lk1 = -7.07277513492202e-8
+ k2 = 0.0227753222192018 lk2 = 2.03511478301116e-08 wk2 = 2.56031459940945e-09 pk2 = -2.9529541923447e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 273386.395625 lvsat = -0.580431349597031
+ ua = 2.61616633625946e-09 lua = 1.36539337636142e-15 wua = -8.29719828904729e-16 pua = 3.23051128841093e-21
+ ub = -1.49686077833208e-19 lub = -1.01584551629779e-24 wub = 9.21918968069361e-25 pub = -5.42586022205092e-30
+ uc = -5.15756313125e-11 luc = 9.17760209583907e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0210016404217217 lu0 = 4.98371762185074e-09 wu0 = -6.0997266816289e-09 pu0 = 4.14821117893795e-15
+ a0 = 0.201965995986916 la0 = 2.64492168679594e-06 wa0 = 3.54899014938349e-06 pa0 = -1.3879937491409e-11
+ keta = -0.00495672689375 lketa = -2.34839323906078e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0383070146285059 lags = 4.49086778523245e-07 wags = 3.87327282050819e-07 pags = -1.55080159715774e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.094776478466875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.24319289368812e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.00300994419849+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.9111312102246e-06 wnfactor = -3.18870488214093e-06 pnfactor = 1.06308639592646e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.64831926658375 lpclm = 5.78838869829003e-06 wpclm = -2.11758236813575e-22 ppclm = -1.61558713389263e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00455412315405625 lpdiblc2 = -1.27602734399944e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 562123300.169375 lpscbe1 = -1806.55551118713
+ pscbe2 = -1.5317388699625e-08 lpscbe2 = 2.39795383634009e-13 ppscbe2 = 9.62964972193618e-35
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.815322348125e-05 lalpha0 = -2.17393918220827e-10
+ alpha1 = 0.0
+ beta0 = 39.1402881918125 lbeta0 = -6.9146000555929e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.53833566097963e-08 lagidl = -8.05273567643065e-14 wagidl = -4.91341360879304e-14 pagidl = 1.63731325650331e-19
+ bgidl = 1342303983.05494 lbgidl = 2030.83980424248 wbgidl = 1039.17276205498 pbgidl = -0.00406238612006343
+ cgidl = 1332.28625 lcgidl = -0.0026281350228125 wcgidl = -1.73472347597681e-18
+ egidl = 1.20931880529937 legidl = -4.07967463450158e-06 wegidl = -1.6940658945086e-21 pegidl = -6.46234853557053e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.879030981290117 lkt1 = 8.19805885641145e-07 wkt1 = -4.09946200961957e-07 pkt1 = -1.59520176094885e-12
+ kt2 = -0.019032
+ at = 648283.313231997 lat = -1.57776339518018 wat = 0.0436942698403735 pat = -3.45588903734975e-7
+ ute = -1.51655375 lute = -1.545961778125e-7
+ ua1 = 2.2096e-11
+ ub1 = -3.27481451126419e-18 lub1 = -3.06788330178373e-24 wub1 = -8.89800528206285e-25 pub1 = 7.03765482771553e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.43 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.864173818371155+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -3.23763587304957e-07 wvth0 = -1.46763415742756e-07 pvth0 = 8.46693854783254e-13
+ k1 = 0.602594105 lk1 = -6.46359499712504e-8
+ k2 = 0.0284159277267564 lk2 = -1.69938925029652e-09 wk2 = -9.06712026569618e-09 pk2 = 1.59250078229671e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 137871.16318875 lvsat = -0.0506684271956208 wvsat = -0.0706621582218883 pvsat = 2.76236042028917e-7
+ ua = 3.32105560571619e-09 lua = -1.39019500026228e-15 wua = -2.03649793394932e-17 pua = 6.65408427480938e-23
+ ub = -1.44260028787921e-18 lub = 4.03847935932453e-24 wub = -6.20778360187988e-25 pub = 6.0492930843913e-31
+ uc = -5.4923007875e-11 luc = 1.04861752785344e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0212519674608157 lu0 = 4.00512664427268e-09 wu0 = -4.37847368333717e-09 pu0 = -2.58059710463412e-15
+ a0 = 0.838751943621997 la0 = 1.55566221003499e-07 wa0 = -3.07066940572547e-08 pa0 = 1.13992393811779e-13
+ keta = -0.00508732849999999 lketa = -2.2973378061375e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.110897808348917 lags = 1.65311218171727e-07 wags = 2.0719596247088e-09 pags = -4.47422279634664e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.064087020519875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.07540834542429e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.57188437596526+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -4.22575358260888e-06 wnfactor = -4.45923098149456e-06 pnfactor = 1.55976681131628e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.019094925 leta0 = 2.3809316444375e-7
+ etab = -0.1224012755 letab = 2.04849686248375e-7
+ dsub = 0.81474168125 ldsub = -9.95848917426563e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04876453907784 lpclm = -8.4593616899256e-07 wpclm = 5.79429697446362e-12 ppclm = -2.26513554470595e-17
+ pdiblc1 = 0.581562116725 lpdiblc1 = -7.48864204807206e-7
+ pdiblc2 = -0.001133342292 lpdiblc2 = 9.473450855001e-9
+ pdiblcb = 0.165925 lpdiblcb = -7.4637355625e-07 wpdiblcb = 5.29395592033938e-23 ppdiblcb = 4.03896783473158e-28
+ drout = 0.139965 ldrout = 1.64202182375e-6
+ pscbe1 = -156170353.9325 lpscbe1 = 1001.43395611063
+ pscbe2 = 7.6074691134375e-08 lpscbe2 = -1.17479104457055e-13
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.4063189874125e-05 lalpha0 = -8.41274543421732e-11
+ alpha1 = -9.54625e-11 lalpha1 = 3.73186778125e-16
+ beta0 = 70.183410779125 lbeta0 = -0.000128269927030044
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.03417799295774e-08 lagidl = -2.17260731271606e-14 wagidl = -3.09532906386571e-14 pagidl = 9.26578555777597e-20
+ bgidl = 2474382862.5 lbgidl = -2394.73955522813
+ cgidl = 842.76295625 lcgidl = -0.000714466086720313
+ egidl = -1.5853225474425 legidl = 6.84527707370459e-06 wegidl = 8.470329472543e-22
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.389566763392364 lkt1 = -1.09363210817565e-06 wkt1 = -3.35929125509577e-06 pkt1 = 9.93452539192377e-12
+ kt2 = -0.019032
+ at = 473279.535420809 lat = -0.893629876771786 wat = -0.560330364659846 pat = 2.01569439868501e-6
+ ute = -1.6575766375 lute = 3.96697545146875e-7
+ ua1 = -4.84145456e-10 lua1 = 1.979024411868e-15 wua1 = 1.97215226305253e-31 pua1 = -9.4039548065783e-37
+ ub1 = -5.26100655978736e-18 lub1 = 4.69663796390549e-24 wub1 = 5.53105503641261e-24 pub1 = -1.80630747882709e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.10187467607197+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.30066775260313e-07 wvth0 = 4.63289405069696e-07 pvth0 = -3.18049493352919e-13
+ k1 = 0.5590564875 lk1 = 1.8488246240625e-8
+ k2 = 0.0261058180026611 lk2 = 2.71118774043248e-09 wk2 = -9.43172623948894e-09 pk2 = 1.66211317784307e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 169019.0178725 lvsat = -0.110137468750571 wvsat = 0.141324316443777 pvsat = -1.28499134726504e-7
+ ua = 3.44848752764965e-09 lua = -1.63349439721373e-15 wua = 3.65244198624953e-17 pua = -4.20752426782995e-23
+ ub = -2.61028670689522e-19 lub = 1.78256374920512e-24 wub = 2.3123975581343e-24 pub = -4.9952368136177e-30
+ uc = 5.32329505e-13 luc = -1.01635010742125e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.025273770378849 lu0 = -3.67350057698244e-09 wu0 = 9.15124635472259e-11 pu0 = -1.11149181555732e-14
+ a0 = 1.02693385851797 la0 = -2.03720100011639e-07 wa0 = -6.22565840579306e-08 pa0 = 1.74229021295567e-13
+ keta = 0.044301656 lketa = -1.17269296718e-07 pketa = -5.04870979341448e-29
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.329814866218907 lags = 1.00674189209035e-06 wags = 1.61729172223986e-07 pags = -3.49567761118636e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.121865847693686+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 2.77339123917048e-09 wvoff = -1.11084363947149e-07 pvoff = 2.12087821866095e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '1.19614290858155+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 2.21938081399348e-06 wnfactor = 9.72917663019554e-06 pnfactor = -1.14915491194565e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.454625e-05 lcit = -8.6799278125e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.285229163291639 leta0 = -2.70023630014561e-07 weta0 = -5.55146548576375e-08 peta0 = 1.05991354786944e-13
+ etab = -0.028844949 letab = 2.622726987825e-8
+ dsub = 0.287839303643931 ldsub = 1.01394470178245e-08 wdsub = 3.36517309735418e-12 pdsub = -6.4249567358621e-18
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0624874866168126 lpclm = 1.03711329341866e-06 wpclm = -1.15885939489272e-11 ppclm = 1.05369290483002e-17
+ pdiblc1 = -0.00178611264999995 lpdiblc1 = 3.64893402127013e-7
+ pdiblc2 = 0.005940118645525 lpdiblc2 = -4.03155443996861e-09 ppdiblc2 = 6.31088724176809e-30
+ pdiblcb = -0.40685 lpdiblcb = 3.471971125e-7
+ drout = 1.5358306539575 ldrout = -1.02303467606836e-06 pdrout = 1.61558713389263e-27
+ pscbe1 = 430963245.09 lpscbe1 = -119.550867823083
+ pscbe2 = 1.4532757728e-08 lpscbe2 = 1.98318990659932e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.165892571425e-05 lalpha0 = 1.17722494844932e-10 walpha0 = -6.37024902488598e-27 palpha0 = 1.86252848108128e-32
+ alpha1 = 1.90925e-10 lalpha1 = -1.7359855625e-16
+ beta0 = -39.87379705625 lbeta0 = 8.18567970296453e-05 pbeta0 = 1.29246970711411e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -4.26601675909514e-09 lagidl = 6.16386270068749e-15 wagidl = 3.33980840826061e-14 pagidl = -3.02050066088121e-20
+ bgidl = 907590775.0 lbgidl = 596.658237831251
+ cgidl = 1306.672187538 lcgidl = -0.00160018478655693 wcgidl = -0.00371515109959567 pcgidl = 7.09315223690303e-9
+ egidl = 3.11021319877 legidl = -2.11967454975162e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.36283133856841 lkt1 = 7.6457328197921e-07 wkt1 = 3.91215473367436e-06 pkt1 = -3.9484828621356e-12
+ kt2 = -0.019032
+ at = -17298.4237696073 lat = 0.0430060918125156 wat = 0.945883649958198 pat = -8.60044708724492e-7
+ ute = -1.43979825 lute = -1.90958411875009e-8
+ ua1 = 5.524e-10
+ ub1 = -2.08291298536853e-18 lub1 = -1.37113719305367e-24 wub1 = -7.50290796000011e-24 pub1 = 6.8220190626301e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.45 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.1511367585406+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.74858323744923e-07 wvth0 = 5.15981991033516e-07 pvth0 = -3.65960227140525e-13
+ k1 = 0.590241525 lk1 = -9.86674910625021e-9
+ k2 = 0.00468799379676071 lk2 = 2.21853443996475e-08 wk2 = 4.02266734758774e-08 pk2 = -2.8530768162766e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9128.48749999993 lvsat = 0.0352429959906251
+ ua = -8.31844341241457e-10 lua = 2.2583973545755e-15 wua = -4.43270695916708e-17 pua = 3.14389741078926e-23
+ ub = 8.47490783940337e-18 lub = -6.16058652259684e-24 wub = -1.44634466694204e-23 pub = 1.02581995502864e-29
+ uc = 6.082695725e-12 luc = -6.06302059295625e-18 wuc = -3.08148791101958e-33 puc = 2.93873587705572e-39
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0297663538249301 lu0 = -7.75838207533169e-09 wu0 = -5.51585522404641e-08 pu0 = 3.91212031765492e-14
+ a0 = 0.658800216729128 la0 = 1.31005413784866e-07 wa0 = 5.88111111204474e-07 pa0 = -4.17117805621772e-13
+ keta = -0.1537600425 lketa = 6.2818302643125e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.977016824904027 lags = -1.8149482306318e-07 wags = -1.01257755636988e-06 pags = 7.18170631855338e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.281923008822819+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.48305364995834e-07 wvoff = 5.55421819735747e-07 pvoff = -3.93932925647578e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.22853720560629+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.44707370057627e-06 wnfactor = -1.32264763422561e-05 pnfactor = 9.38087834574516e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.273125e-05 lcit = 1.61221390625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0559184715706923 leta0 = 4.01648569840135e-08 weta0 = 2.77573274288187e-07 peta0 = -1.96868844788897e-13
+ etab = 0.0018863213 letab = -1.715137642025e-9
+ dsub = 0.384693796942844 ldsub = -7.79255010142126e-08 wdsub = -1.68258654859239e-11 pdsub = 1.19337450960291e-17
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.0219588243125 lpclm = -7.4453602038114e-7
+ pdiblc1 = 0.1958620354125 lpdiblc1 = 1.85181823501184e-7
+ pdiblc2 = -0.033618504135125 lpdiblc2 = 3.19371233233374e-08 wpdiblc2 = -1.98523347012727e-23 ppdiblc2 = 6.31088724176809e-30
+ pdiblcb = -0.025
+ drout = 0.335842470275 ldrout = 6.80545799449562e-8
+ pscbe1 = -56987686.1249995 lpscbe1 = 324.118516384156
+ pscbe2 = 1.82815146225e-08 lpscbe2 = -3.38872530725814e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0002471576267875 lalpha0 = -1.63068955517284e-10 palpha0 = 1.97215226305253e-31
+ alpha1 = 0.0
+ beta0 = 67.19689401875 lbeta0 = -1.54972288302985e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.91011851875989e-08 lagidl = 1.96527395943045e-14 wagidl = 8.11006716487821e-16 pagidl = -5.75206513668999e-22
+ bgidl = 700288124.999998 lbgidl = 785.148172343748
+ cgidl = -3904.51550018999 lcgidl = 0.00313808761850975 wcgidl = 0.0185757554979783 pcgidl = -1.31748545869411e-8
+ egidl = 1.8355566512875 legidl = -9.6069308395316e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.70546585057057 lkt1 = 1.07611371201717e-06 wkt1 = -1.95678085271095e-06 pkt1 = 1.38784681978524e-12
+ kt2 = -0.019032
+ at = 47731.25 lat = -0.0161221390625
+ ute = -1.39342125 lute = -6.12641284375002e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.46 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.497079867157968+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.89031526468211e-07 wvth0 = -1.18977107733753e-06 pvth0 = 8.43845136601641e-13
+ k1 = 0.621240645643238 lk1 = -3.18528754224665e-08 wk1 = -1.33629200936589e-07 pk1 = 9.47765107642751e-14
+ k2 = 0.0253229954909538 lk2 = 7.54996944804107e-09 wk2 = -2.45018280983856e-10 pk2 = 1.73779215787835e-16
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 119228.373515168 lvsat = -0.0428453481656329 wvsat = -0.292316232993797 pvsat = 2.0732528825085e-7
+ ua = -8.55857795844092e-09 lua = 7.73858317257422e-15 wua = 3.2524201576313e-14 pua = -2.3067789968e-20
+ ub = 5.75923497954808e-18 lub = -4.23449554674448e-24 wub = -1.67840424998204e-23 pub = 1.19040821429976e-29
+ uc = 1.05905924964515e-11 luc = -9.26024637810822e-18 wuc = -3.88485908279966e-17 puc = 2.75533630447566e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.0200170832193702 lu0 = 2.75505206483383e-08 wu0 = 1.25264653775001e-07 pu0 = -8.88439556899191e-14
+ a0 = 1.08123870676879 la0 = -1.68609085275762e-07 wa0 = -7.07348929640361e-07 pa0 = 5.01687228347426e-13
+ keta = 0.21966793817985 lketa = -2.02035492654058e-07 wketa = -1.01550653687777e-06 pketa = 7.20248011280558e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -2.6289987965861 lags = 2.37607175647869e-06 wags = 9.96809757282692e-06 pags = -7.06987320352749e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '0.13650667525959+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.48465888439614e-07 wvoff = -6.22844178913073e-07 pvoff = 4.41752233894096e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.95406600452658+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.96165500121047e-06 wnfactor = -5.01835134575121e-06 pnfactor = 3.55926569197405e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.146754257435802 leta0 = 1.04590138108842e-07 weta0 = 4.42334706745396e-07 peta0 = -3.13725890759172e-13
+ etab = -0.0018863213 letab = 9.60609122025e-10
+ dsub = 0.0621317022650203 ldsub = 1.50851664636034e-07 wdsub = 6.32879581122931e-07 pdsub = -4.48869842911437e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.894842824149528 lpclm = 1.32420554879055e-06 wpclm = 5.55529006096728e-06 ppclm = -3.94008947574104e-12
+ pdiblc1 = -0.241109631949019 lpdiblc1 = 4.95103978577341e-07 wpdiblc1 = 2.07706049015444e-06 ppdiblc1 = -1.47315515264204e-12
+ pdiblc2 = 0.0494858065169306 lpdiblc2 = -2.70046090066331e-08 wpdiblc2 = -1.13289750934579e-07 ppdiblc2 = 8.03507558503504e-14
+ pdiblcb = -0.025
+ drout = -2.4791387589403 ldrout = 2.06458001676591e-06 wdrout = 8.66132725070998e-06 pdrout = -6.14304635256605e-12
+ pscbe1 = 480165439.129532 lpscbe1 = -56.8573377026207 wpscbe1 = -238.527935196209 ppscbe1 = 0.000169175938037912
+ pscbe2 = 6.14496453798506e-09 lpscbe2 = 5.2191228401841e-15 wpscbe2 = 2.18952670826005e-14 ppscbe2 = -1.55292181783344e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000328250996553267 lalpha0 = 2.45039610587154e-10 walpha0 = 1.0279903125317e-09 palpha0 = -7.29102129163107e-16
+ alpha1 = 0.0
+ beta0 = -1.62343297194951 lbeta0 = 3.33135880878552e-05 wbeta0 = 0.000139757183534235 pbeta0 = -9.91227824216565e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.73702413117569e-08 lagidl = -6.21461965036356e-15 wagidl = -9.19779779253378e-15 pagidl = 6.52353808435459e-21
+ bgidl = 2441369905.34387 lbgidl = -449.714080365143 wbgidl = -1886.64076357581 pbgidl = 0.00133809996156614
+ cgidl = 2356.9657597375 lcgidl = -0.00130286796509382 wcgidl = -0.0054657924219479 pcgidl = 3.87661327526655e-9
+ egidl = -1.32948408403491 legidl = 1.28411205757426e-06 wegidl = 5.38710762814394e-06 pegidl = -3.82080608526109e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 1.76639686103176 lkt1 = -1.38630491618678e-06 wkt1 = -5.25207993824974e-06 pkt1 = 3.72503769620363e-12
+ kt2 = -0.019032
+ at = 42823.75 lat = -0.0126414946875
+ ute = -1.7271215656625 lute = 1.75412820446128e-07 wute = 5.65426802270479e-07 pute = -4.01028959510332e-13
+ ua1 = 5.53418499999999e-10 lua1 = -7.22371125000165e-19
+ ub1 = -4.333641125e-18 lub1 = 5.26789142906246e-25
+ uc1 = -2.8159131e-10 luc1 = 1.222685366175e-16 puc1 = 1.88079096131566e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.47 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.184632154569+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 6.11044758958572e-08 wvth0 = 1.78049739344485e-06 pvth0 = -6.68764082144284e-13
+ k1 = 0.338079641278201 lk1 = 1.12346866050429e-07 wk1 = 8.01324603667796e-07 pk1 = -3.81348714230505e-13
+ k2 = 0.0746133794655651 lk2 = -1.75511585910297e-08 wk2 = -1.37010047949988e-07 pk2 = 6.98213705747279e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 226088.529144955 lvsat = -0.0972638824201018 wvsat = -1.06017026340102 pvsat = 5.9835495323573e-7
+ ua = 2.08376954887961e-08 lua = -7.23146908043124e-15 wua = -5.81859762921062e-14 pua = 2.31263681114925e-20
+ ub = -1.49549885966426e-17 lub = 6.31422280943061e-24 wub = 3.63114222222454e-23 pub = -1.51347832667144e-29
+ uc = -1.57596604579196e-10 luc = 7.63890837326654e-17 wuc = 8.69929713090672e-16 puc = -4.35241988225826e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0700208335919499 lu0 = -1.83012884878265e-08 wu0 = -1.85255996886761e-07 pu0 = 6.92886856595831e-14
+ a0 = 1.3237196009585 la0 = -2.92092480641874e-07 wa0 = -2.43039703543231e-06 pa0 = 1.37914947622198e-12
+ keta = -0.137049892726472 lketa = -2.03769372650138e-08 wketa = -2.33178007247698e-07 pketa = 3.21847207566444e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.1969005669778 lags = 1.64677573305067e-06 wags = 1.21744216383674e-05 pags = -8.193443733904e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.169010859916058+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 7.11891634858414e-09 wvoff = 8.65734031982967e-07 pvoff = -3.16306220004712e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '0.916622653758747+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 6.03663025168042e-07 wnfactor = 1.34670859411463e-05 pnfactor = -5.85444324637853e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 6.09050318875e-05 lcit = -2.59233874887094e-11 wcit = -1.51465173509534e-10 pcit = 7.71336396097304e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.763513097995662 leta0 = -3.5896351264463e-07 weta0 = -4.0191805932012e-06 peta0 = 1.95830077573863e-12
+ etab = 0.0121563598841775 letab = -6.19062627101742e-09 wetab = 1.47799716310604e-07 petab = -7.52670055311749e-14
+ dsub = 0.652297114065168 ldsub = -1.49690071323191e-07 wdsub = -1.3463674129359e-06 pdsub = 5.5906168881302e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.316549529527554 lpclm = 7.07303992680498e-07 wpclm = 6.41400103918796e-06 ppclm = -4.37738804139993e-12
+ pdiblc1 = 0.877940138667317 lpdiblc1 = -7.47721171090276e-08 wpdiblc1 = 2.00625783359632e-06 ppdiblc1 = -1.43709889978981e-12
+ pdiblc2 = -0.0758644600276356 lpdiblc2 = 3.68300142311873e-08 wpdiblc2 = 3.52014155413871e-07 ppdiblc2 = -1.56605258457598e-13
+ pdiblcb = -1.2427012755 lpdiblcb = 6.20114374548375e-07 wpdiblcb = 6.05860694038137e-06 ppdiblcb = -3.08534558438921e-12
+ drout = 6.75183483059918 ldrout = -2.63629328370707e-06 wdrout = -2.57239714628912e-05 pdrout = 1.13676670173354e-11
+ pscbe1 = 886035991.106242 lpscbe1 = -263.54691629676 wpscbe1 = -1060.72974651373 ppscbe1 = 0.000587882210451359
+ pscbe2 = 2.48209480061787e-08 lpscbe2 = -4.2916217409935e-15 wpscbe2 = -4.63324832931074e-14 ppscbe2 = 1.92157637004949e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000329985245720384 lalpha0 = -9.01671957907021e-11 walpha0 = -7.20623517132361e-10 palpha0 = 1.61379463593315e-16
+ alpha1 = 6.0885063775e-10 lalpha1 = -3.10057187274188e-16 walpha1 = -3.02930347019069e-15 palpha1 = 1.54267279219461e-21
+ beta0 = -171.353305738435 lbeta0 = 0.000119748525794188 wbeta0 = 0.00116043592588032 pbeta0 = -6.18903431961402e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.80462707745982e-08 lagidl = -1.67438876543155e-14 wagidl = -2.08977258419811e-13 pagidl = 1.08261228408795e-19
+ bgidl = -1656484391.4045 lbgidl = 1637.11822025397 wbgidl = 17456.645302003 pbgidl = -0.00851246846732984
+ cgidl = -419.70399987645 lcgidl = 0.000111151109989582 wcgidl = -0.000228975000980717 pcgidl = 1.20976400363901e-9
+ egidl = 11.3823929755749 legidl = -5.18941133503202e-06 wegidl = -5.09328283120472e-05 pegidl = 2.48601212922812e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -2.46453326801357 lkt1 = 7.68296252029557e-07 wkt1 = 9.87454944325505e-06 pkt1 = -3.97819831632769e-12
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -0.815840730924997 lute = -2.88656944643944e-07 wute = -4.16015707473163e-06 pute = 2.00547462985299e-12
+ ua1 = 5.52e-10
+ ub1 = -4.957481e-18 lub1 = 8.44479599250001e-25
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.48 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.90589393478+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = -1.78677472885882e-8
+ k1 = 0.608803775813334 wk1 = -4.04475458686794e-8
+ k2 = 0.0241669092301427 wk2 = 2.34224362740893e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 219328.3426 wvsat = -0.0575104396757996
+ ua = 2.61614232689791e-09 wua = 9.24574412477322e-17
+ ub = -2.02302379946667e-19 wub = 1.03021245627897e-26
+ uc = -5.60297706333333e-11 wuc = 4.77790293998691e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0199184301617333 wu0 = -4.7735128300881e-10
+ a0 = 1.31601157621213 wa0 = -5.25676734754087e-7
+ keta = -0.00625884274613333 wketa = -4.96023883778856e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.169665996769493 wags = -3.06530350798018e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0874903097253173+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' wvoff = -1.70027317410655e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.19125460053333+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = -1.65302271393851e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.49181533333333e-05 wcit = -1.46336996630533e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.66221915003436 wpclm = 2.21894004478064e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00456455310587613 wpdiblc2 = -4.83142628185252e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 447221920.362453 wpscbe1 = -337.740168882601
+ pscbe2 = 1.501649444638e-08 wpscbe2 = -4.62278572355832e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.06839939075347e-05 walpha0 = -8.93133820949044e-11
+ alpha1 = 0.0
+ beta0 = 39.0497950461547 wbeta0 = -2.33200296438472e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.46198057373333e-09 wagidl = -5.40305458959255e-15
+ bgidl = 1758978278.66667 wbgidl = 49.7545788543812
+ cgidl = 1523.29151466667 wcgidl = -0.00155702564414887
+ egidl = 0.49835708641752 wegidl = 5.80661749076835e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.11357275909333 wkt1 = 3.94641612513222e-7
+ kt2 = -0.019032
+ at = 554274.716386667 wat = -0.313834322973842
+ ute = -1.51642738666667 wute = -5.85347986522143e-8
+ ua1 = 2.2096e-11
+ ub1 = -3.5732879724e-18 wub1 = -2.66040659874311e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.49 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.90589393478+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = -1.78677472885886e-8
+ k1 = 0.608803775813333 wk1 = -4.04475458686798e-8
+ k2 = 0.0241669092301427 wk2 = 2.34224362740891e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 219328.3426 wvsat = -0.0575104396757995
+ ua = 2.61614232689791e-09 wua = 9.24574412477322e-17
+ ub = -2.02302379946667e-19 wub = 1.03021245627896e-26
+ uc = -5.60297706333333e-11 wuc = 4.77790293998691e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0199184301617333 wu0 = -4.77351283008796e-10
+ a0 = 1.31601157621213 wa0 = -5.25676734754088e-7
+ keta = -0.00625884274613333 wketa = -4.96023883778855e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.169665996769493 wags = -3.06530350798018e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0874903097253173+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' wvoff = -1.70027317410654e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.19125460053333+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = -1.6530227139385e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.49181533333333e-05 wcit = -1.46336996630533e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.66221915003436 wpclm = 2.21894004478064e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00456455310587613 wpdiblc2 = -4.83142628185252e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 447221920.362453 wpscbe1 = -337.7401688826
+ pscbe2 = 1.501649444638e-08 wpscbe2 = -4.62278572355832e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.06839939075347e-05 walpha0 = -8.93133820949044e-11
+ alpha1 = 0.0
+ beta0 = 39.0497950461547 wbeta0 = -2.33200296438472e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.46198057373333e-09 wagidl = -5.40305458959255e-15
+ bgidl = 1758978278.66667 wbgidl = 49.7545788543812
+ cgidl = 1523.29151466667 wcgidl = -0.00155702564414887
+ egidl = 0.49835708641752 wegidl = 5.80661749076836e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.11357275909333 wkt1 = 3.94641612513223e-7
+ kt2 = -0.019032
+ at = 554274.716386667 wat = -0.313834322973842
+ ute = -1.51642738666667 wute = -5.85347986522134e-8
+ ua1 = 2.2096e-11
+ ub1 = -3.5732879724e-18 wub1 = -2.66040659874311e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.50 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.883351579490081+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.78293123576792e-07 wvth0 = -5.11277752316778e-08 pvth0 = 2.63061876008884e-13
+ k1 = 0.626542213283471 lk1 = -1.40297736560685e-07 wk1 = -6.6619652480244e-08 pk1 = 2.07001734217516e-13
+ k2 = 0.0215518952079057 lk2 = 2.06827996553779e-08 wk2 = 6.20055560646243e-09 pk2 = -3.05163540203288e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 364899.847477883 lvsat = -1.15136142495539 wvsat = -0.272293334261852 pvsat = 1.69877160900473e-6
+ ua = 2.00140510583548e-09 lua = 4.86211036568804e-15 wua = 9.99469015115411e-16 pua = -7.17378129061295e-21
+ ub = 5.09813492829903e-19 lub = -5.63230246675808e-24 wub = -1.04038639146191e-24 pub = 8.31015814536835e-30
+ uc = -7.90470895495019e-11 luc = 1.82049729637707e-16 wuc = 8.17398405254544e-17 puc = -2.68604545395036e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0183188689861475 lu0 = 1.26513292280023e-08 wu0 = 1.88271485526464e-09 pu0 = -1.86663531041391e-14
+ a0 = 1.82260118863798 la0 = -4.00674389207915e-06 wa0 = -1.27312235204936e-06 pa0 = 5.91173424859262e-12
+ keta = -0.000369099917933904 lketa = -4.65834484639364e-08 wketa = -1.36502363346841e-08 pketa = 6.8731362702321e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.187751836206259 lags = -1.4304542556524e-07 wags = -5.73377145334202e-08 pags = 2.11055800968531e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0906082229895355+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 2.46603554850181e-08 wvoff = -1.24024190870276e-08 pvoff = -3.6385022858948e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.77768928192312+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -4.63825850378221e-06 wnfactor = -2.51827541885635e-06 pnfactor = 6.84349995637145e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.49181533333333e-05 wcit = -1.46336996630533e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.11394027814573 lpclm = 1.14820253325148e-05 wpclm = 4.36087617636805e-06 ppclm = -1.69411083487577e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00776481478816271 lpdiblc2 = -2.53116697106251e-08 wpdiblc2 = -9.55323957993551e-09 ppdiblc2 = 3.73460018278629e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 900303933.578178 lpscbe1 = -3583.53891302647 wpscbe1 = -1006.23821295369 ppscbe1 = 0.00528731815506925
+ pscbe2 = -4.51239078296283e-08 lpscbe2 = 4.75665476701519e-13 wpscbe2 = 8.86876881192918e-14 ppscbe2 = -7.01818724937349e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0001352061348096 lalpha0 = -4.31229242929657e-10 walpha0 = -1.69757856800293e-10 palpha0 = 6.36255461563591e-16
+ alpha1 = 0.0
+ beta0 = 40.7839686679278 lbeta0 = -1.37160127180094e-05 wbeta0 = -4.89068249793543e-06 pbeta0 = 2.0237236100736e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.38573173355078e-08 lagidl = -5.05823172830649e-14 wagidl = -1.48390286334057e-14 pagidl = 7.4631477706029e-20
+ bgidl = 1592062490.01324 lbgidl = 1320.1787014071 wbgidl = 296.029811559925 pbgidl = -0.0019478523842763
+ cgidl = 2182.42471027833 lcgidl = -0.00521324922739158 wcgidl = -0.00252954108108133 pcgidl = 7.691867719558e-9
+ egidl = 1.52153472209972 legidl = -8.09256771501947e-06 wegidl = -9.28981600779929e-07 pegidl = 1.19401466648546e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.18472037167848 lkt1 = 5.62724254839033e-07 wkt1 = 4.99616072911519e-07 pkt1 = -8.30269250905233e-13
+ kt2 = -0.019032
+ at = 979105.447228845 lat = -3.3600924579135 wat = -0.940649125472011 pat = 4.95763497665864e-6
+ ute = -1.47765484574833 lute = -3.0666171925833e-07 wute = -1.15741589060005e-07 pute = 4.52462807032821e-13
+ ua1 = 2.2096e-11
+ ub1 = -3.39706677392617e-18 lub1 = -1.3937775140291e-24 wub1 = -5.26045522277721e-25 pub1 = 2.05644345796418e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.51 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.911056815753552+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -6.99864287138172e-08 wvth0 = -7.26558871329155e-09 pvth0 = 9.15936233618832e-14
+ k1 = 0.62345111293722 lk1 = -1.28213852532104e-07 wk1 = -6.20589008387703e-08 pk1 = 1.89172615863083e-13
+ k2 = 0.0229891772820937 lk2 = 1.50641047068583e-08 wk2 = 7.07988263787368e-09 pk2 = -3.39538632178732e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 48979.5711356166 lvsat = 0.0836499153356105 wvsat = 0.193829973786239 pvsat = -1.23420932982265e-7
+ ua = 3.93891150214322e-09 lua = -2.71208651407802e-15 wua = -1.85876183493972e-15 pua = 3.99975765996508e-21
+ ub = -3.00720984673159e-18 lub = 8.11662102342269e-24 wub = 4.0346328932611e-24 pub = -1.15293609934351e-29
+ uc = -9.78301759860135e-11 luc = 2.55477510289639e-16 wuc = 1.27667961727243e-16 puc = -4.48149053203126e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0201009413649824 lu0 = 5.68476278104206e-09 wu0 = -9.5365769059427e-10 pu0 = -7.57826372924023e-15
+ a0 = 0.605351771014418 la0 = 7.51788393765771e-07 wa0 = 6.63762915927274e-07 pa0 = -1.66003448524503e-12
+ keta = -0.00062816526920733 lketa = -4.55706972394707e-08 wketa = -1.32679993984091e-08 pketa = 6.72371029591881e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0758409515231108 lags = 2.94442200382358e-07 wags = 1.06381744039628e-07 pags = -4.28964492458157e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0297316730624893+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -2.13321297317288e-07 wvoff = -1.02222481170688e-07 pvoff = 3.14744054841603e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.88580030213886+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 2.75760849043943e-06 wnfactor = 5.5762113163593e-07 pnfactor = -5.18094863364049e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.49181533333333e-05 wcit = -1.46336996630533e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0408131745256334 leta0 = 4.72288902514333e-07 weta0 = 1.78253315101148e-07 peta0 = -6.96836772059162e-13
+ etab = -0.173944777054249 letab = 4.06346119699322e-07 wetab = 1.53364905525583e-07 petab = -5.99541756925886e-13
+ dsub = 1.06531341100573 ldsub = -1.97539645197413e-06 wdsub = -7.45562651014753e-07 pdsub = 2.91459079347943e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.25245106553263 lpclm = -1.67804002775979e-06 wpclm = -6.06052466096819e-07 ppclm = 2.47585744679807e-12
+ pdiblc1 = 0.76998848930729 lpdiblc1 = -1.48547000182452e-06 wpdiblc1 = -5.60652496594484e-07 ppdiblc1 = 2.19173077231199e-12
+ pdiblc2 = -0.00351701608624149 lpdiblc2 = 1.87918276351396e-08 wpdiblc2 = 7.09249265638066e-09 ppdiblc2 = -2.77263269169561e-14
+ pdiblcb = 0.353724685033333 lpdiblcb = -1.48052947496656e-06 wpdiblcb = -5.58787821633692e-07 ppdiblcb = 2.18444129172151e-12
+ drout = -0.273194307073333 ldrout = 3.25716484492643e-06 wdrout = 1.22933320759412e-06 pdrout = -4.80577084178732e-12
+ pscbe1 = -524525386.370361 lpscbe1 = 1986.47510598236 wpscbe1 = 1096.0205078471 ppscbe1 = -0.00293093674922125
+ pscbe2 = 1.36164224419542e-07 lpscbe2 = -2.33035154293552e-13 wpscbe2 = -1.78793161455218e-13 ppscbe2 = 3.43830786261804e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.75840987188092e-05 lalpha0 = -1.66877798341735e-10 walpha0 = -6.99851941382801e-11 palpha0 = 2.46219180052119e-16
+ alpha1 = -1.89362342516667e-10 lalpha1 = 7.4026473748328e-16 walpha1 = 2.79393910816846e-16 palpha1 = -1.09222064586076e-21
+ beta0 = 102.362058621214 lbeta0 = -0.000254440160867892 wbeta0 = -9.57458290071512e-05 pbeta0 = 3.75412717591888e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.59395283237199e-10 lagidl = 2.57535949977404e-15 wagidl = -9.53699572242695e-16 pagidl = 2.03502550736776e-20
+ bgidl = 2964713233.20663 lbgidl = -4045.85621642167 wbgidl = -1458.95154019757 pbgidl = 0.00491280846508168
+ cgidl = 1898.73813997016 lcgidl = -0.00410424750241435 wcgidl = -0.00314199713649941 pcgidl = 1.00861115542011e-8
+ egidl = -4.02200156753388 legidl = 1.35785015252307e-05 wegidl = 7.25020684361481e-06 pegidl = -2.00343457613955e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -2.15132899305234 lkt1 = 4.34143900794483e-06 wkt1 = 1.88273712409709e-06 pkt1 = -6.23723522025243e-12
+ kt2 = -0.019032
+ at = 182263.845965143 lat = -0.245039428173373 wat = 0.305571104468255 pat = 8.58485427646554e-8
+ ute = -1.62001670049333 lute = 2.49866361403562e-07 wute = -1.11757564326738e-07 pute = 4.36888258344303e-13
+ ua1 = -4.84145456e-10 lua1 = 1.979024411868e-15 wua1 = -4.93038065763132e-32 pua1 = -9.4039548065783e-38
+ ub1 = -3.52520976853935e-18 lub1 = -8.92834512337546e-25 wub1 = 3.66285417080886e-25 pub1 = -1.43190126672345e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.52 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.987352493350997+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 7.56810937391031e-08 wvth0 = 1.22534834581322e-07 pvth0 = -1.5622783481336e-13
+ k1 = 0.537088559710617 lk1 = 3.66738522157884e-08 wk1 = 6.53643828692091e-08 pk1 = -5.41102885563761e-14
+ k2 = 0.0232693516803531 lk2 = 1.45291817369816e-08 wk2 = -9.91973866642734e-10 pk2 = -1.85426711866254e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 225258.741820957 lvsat = -0.252911091295376 wvsat = -0.0260139452197637 pvsat = 2.96316069379946e-7
+ ua = 4.23069980081529e-09 lua = -3.26918332331767e-15 wua = -2.29090595947912e-15 pua = 4.82482882974194e-21
+ ub = 1.15650654101796e-18 lub = 1.67045510111857e-25 wub = -1.90540191739988e-24 pub = -1.88349531180603e-31
+ uc = 6.84425553192915e-11 luc = -6.19787019550142e-17 wuc = -2.0206320975823e-16 puc = 1.81390185955513e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0306362547253528 lu0 = -1.44297842522452e-08 wu0 = -1.58642701353203e-08 pu0 = 2.08898230808529e-14
+ a0 = 1.14854311167707 la0 = -2.85299673394392e-07 wa0 = -4.24098349933151e-07 pa0 = 4.16964636598987e-13
+ keta = 0.0973413389805174 lketa = -2.32618973228258e-07 wketa = -1.57816712565648e-07 pketa = 3.4321673357374e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.705658861627077 lags = 1.78652071863935e-06 wags = 1.28003268498524e-06 pags = -2.66975755145857e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.218399769159928+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.46893265156747e-07 wvoff = 1.76147106543893e-07 pvoff = -2.16733080502461e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.27539528928262+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.80472573876479e-06 wnfactor = -2.40841854895192e-06 pnfactor = 4.81962626521866e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.39362342516667e-05 lcit = -1.72177709933279e-11 wcit = -2.79393910816846e-11 pcit = 2.54038913410217e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.450089092094544 leta0 = -4.64966250030241e-07 weta0 = -5.46046470574526e-07 peta0 = 6.86032593742118e-13
+ etab = 0.0116364212518307 letab = 5.20252168334397e-08 wetab = -1.20450131190329e-07 petab = -7.67603980760312e-14
+ dsub = 0.0201359398954783 ldsub = 2.01086347431075e-08 wdsub = 7.96540268024976e-07 pdsub = -2.96692046971794e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.703971933532877 lpclm = 2.05726058320604e-06 wpclm = 2.28054702725277e-06 ppclm = -3.03538263587963e-12
+ pdiblc1 = -0.387158947826661 lpdiblc1 = 7.23813742523474e-07 wpdiblc1 = 1.14665606093506e-06 ppdiblc1 = -1.06794809115129e-12
+ pdiblc2 = 0.0105141179489019 lpdiblc2 = -7.99711502145789e-09 wpdiblc2 = -1.36096879312354e-08 ppdiblc2 = 1.179931136995e-14
+ pdiblcb = -0.782449370066667 lpdiblcb = 6.88710839733117e-07 wpdiblcb = 1.11757564326738e-06 ppdiblcb = -1.01615565364087e-12
+ drout = 2.49568761066349 ldrout = -2.02932295651259e-06 wdrout = -2.856002542403e-06 pdrout = 2.99415643889468e-12
+ pscbe1 = 640130826.08104 lpscbe1 = -237.14476764048 wpscbe1 = -622.366842189467 ppscbe1 = 0.000349894298836075
+ pscbe2 = 1.40877580286991e-08 lpscbe2 = 3.93391631655581e-17 wpscbe2 = 1.32407257528599e-15 ppscbe2 = -5.80428109359714e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.00014212953190717 lalpha0 = 2.33517950930916e-10 walpha0 = 2.39435943314298e-10 palpha0 = -3.44543126629216e-16
+ alpha1 = 3.78724685033333e-10 lalpha1 = -3.44355419866559e-16 walpha1 = -5.58787821633692e-16 palpha1 = 5.08077826820434e-22
+ beta0 = -115.950793928743 lbeta0 = 0.000162373652863113 wbeta0 = 0.000226362996036273 pbeta0 = -2.39573556622269e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.96447729032663e-10 lagidl = 2.50461711763906e-15 wagidl = 1.98227173712642e-14 pagidl = -1.93171189757129e-20
+ bgidl = 209898641.422866 lbgidl = 1213.77354294149 wbgidl = 2075.94526808355 pbgidl = -0.00183619326612905
+ cgidl = -1623.25367585765 lcgidl = 0.0026201153719549 wcgidl = 0.00500268509094147 pcgidl = -5.46412298854036e-9
+ egidl = 5.29220713508279 legidl = -4.20465144024018e-06 wegidl = -6.49240512982614e-06 pegidl = 6.20373614889661e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.695016479124458 lkt1 = -1.09294608480873e-06 wkt1 = -2.21086032408861e-06 pkt1 = 1.57846570769612e-12
+ kt2 = -0.019032
+ at = 57782.9960622432 lat = -0.00737436549626114 wat = 0.722482939645198 pat = -7.10140378546921e-7
+ ute = -1.45231249115667 lute = -7.03229002724673e-08 wute = 3.72354487926408e-08 pute = 1.52423348046131e-13
+ ua1 = 5.524e-10
+ ub1 = -4.3583154379213e-18 lub1 = 6.97772486929941e-25 wub1 = -7.32570834161766e-25 pub1 = 6.66090030961588e-31
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.53 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.901605942292811+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.2839578105505e-09 wvth0 = -2.2648347804771e-07 pvth0 = 1.61117065944586e-13
+ k1 = 0.583495429321883 lk1 = -5.52159397825579e-09 wk1 = 2.00726434010684e-08 pk1 = -1.292877444497e-14
+ k2 = 0.0398095265908075 lk2 = -5.09972300349095e-10 wk2 = -6.42755507900382e-08 pk2 = 3.8997921130972e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -455963.277341425 lvsat = 0.36649002962802 wvsat = 1.38385543133036 pvsat = -9.85607661248253e-7
+ ua = -8.83979800802908e-09 lua = 8.61516680937407e-15 wua = 2.37829066364369e-14 pua = -1.88827852730947e-20
+ ub = 1.04698980639232e-17 lub = -8.30115573208973e-24 wub = -2.03994323530071e-23 pub = 1.66273476423952e-29
+ uc = 1.20166401209316e-11 luc = -1.06734385609055e-17 wuc = -1.76561311170972e-17 puc = 1.37180497010628e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.00995640817569698 lu0 = 2.24790944905343e-08 wu0 = 6.30343810632536e-08 pu0 = -5.08487755214505e-14
+ a0 = 0.638078905035741 la0 = 1.78839906494234e-07 wa0 = 6.49766255197319e-07 pa0 = -5.59446755615894e-13
+ keta = -0.487378027556905 lketa = 2.99037110795894e-07 wketa = 9.92662299165629e-07 pketa = -7.02856307842924e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 3.21821407722305 lags = -1.78126075101013e-06 wags = -7.68113895599352e-06 pags = 5.47818776310137e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0378417446554652+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.72791186239359e-08 wvoff = -1.70828801405948e-07 pvoff = 9.87547638009314e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '-0.220686133723593+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 3.19258629510361e-06 wnfactor = 2.98739344585962e-06 pnfactor = -4.42417942976052e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.273125e-05 lcit = 1.61221390625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.259815042824538 leta0 = 1.80514084644935e-07 weta0 = 8.84256511639158e-07 peta0 = -6.14470392835674e-13
+ etab = 0.302487493130751 letab = -2.12431120272468e-07 wetab = -8.94422554319119e-07 petab = 6.26974027653822e-13
+ dsub = -0.816055110550594 ldsub = 7.80415347361199e-07 wdsub = 3.57274670794023e-06 pdsub = -2.55393491019013e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.26770631928296 lpclm = -2.46323786816676e-06 wpclm = -6.68210040091986e-06 ppclm = 5.11390453818633e-12
+ pdiblc1 = 0.228614075292368 lpdiblc1 = 1.63922121252497e-07 wpdiblc1 = -9.7451926052393e-08 ppdiblc1 = 6.32570960170468e-14
+ pdiblc2 = -0.0494207478878231 lpdiblc2 = 4.64986617405843e-08 wpdiblc2 = 4.70187229649905e-08 ppdiblc2 = -4.33270712374435e-14
+ pdiblcb = -0.025
+ drout = 0.0668626154906704 ldrout = 1.79086170348289e-07 wdrout = 8.00335032998614e-07 pdrout = -3.30368501539237e-13
+ pscbe1 = 197557456.754715 lpscbe1 = 165.265068419482 wpscbe1 = -757.385327200876 ppscbe1 = 0.0004726598563327
+ pscbe2 = 1.62888022760051e-08 lpscbe2 = -1.96196031869739e-15 wpscbe2 = 5.92920798052892e-15 ppscbe2 = -4.24526217815309e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000513370145671293 lalpha0 = -3.62495130907301e-10 walpha0 = -7.92100974462705e-10 palpha0 = 5.93381815859525e-16
+ alpha1 = 0.0
+ beta0 = 131.244395370038 lbeta0 = -6.23885730068033e-05 wbeta0 = -0.000190569881705684 pbeta0 = 1.39522662464605e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.2055015394748e-08 lagidl = 3.19201849629366e-14 wagidl = 3.93544289910288e-14 pagidl = -3.70763277659839e-20
+ bgidl = 548752443.570002 lbgidl = 905.67072333921 wbgidl = 450.886237168168 pbgidl = -0.000358608342269242
+ cgidl = 3841.92783339 lcgidl = -0.00234910091532852 wcgidl = -0.00447336833314894 pcgidl = 3.15197858731384e-9
+ egidl = 0.218104400613138 legidl = 4.08976471076351e-07 wegidl = 4.81264182946003e-06 pegidl = -4.07537779883434e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -3.29106616762038 lkt1 = 2.53139956174401e-06 wkt1 = 2.76108726825366e-06 pkt1 = -2.94227764064109e-12
+ kt2 = -0.019032
+ at = 119726.867108333 lat = -0.0636968302449187 wat = -0.214219070942522 pat = 1.41555924579963e-7
+ ute = -1.70644941428333 lute = 1.60751097080453e-07 wute = 9.3139839930419e-07 pute = -6.60594314706494e-13
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.54 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.865033521530613+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.822294723614e-08 wvth0 = -9.4944848249058e-08 pvth0 = 6.78232927598932e-14
+ k1 = 0.70191557406815 lk1 = -8.9511081639545e-08 wk1 = -3.7367309401878e-07 pk1 = 2.66335389820058e-13
+ k2 = -0.00363173216900381 lk2 = 3.03007404750472e-08 wk2 = 8.59082103159264e-08 pk2 = -6.75199114334334e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 22554.558733982 lvsat = 0.027101254391538 wvsat = -0.00466851749837571 pvsat = -7.97050541473752e-10
+ ua = 2.89377098995614e-09 lua = 2.9313299755306e-16 wua = -1.55164429279925e-15 pua = -9.14255026533968e-22
+ ub = -5.37428333762268e-19 lub = -4.94209484531315e-25 wub = 1.95133916911565e-24 pub = 7.75062940329696e-31
+ uc = -5.19633150204846e-12 luc = 1.53486156269312e-18 wuc = 8.12454903564408e-18 puc = -4.56689769726899e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0255068275642672 lu0 = -2.67320545803525e-09 wu0 = -1.01892844705302e-08 pu0 = 1.08510925838575e-15
+ a0 = 1.00544265757667 la0 = -8.17128349954172e-08 wa0 = -4.81821878255864e-07 pa0 = 2.43132128035775e-13
+ keta = -0.14481252411372 lketa = 5.60725274788149e-08 wketa = 6.89853967317842e-08 pketa = -4.77384647917201e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.672843756388567 lags = 2.40431490417319e-08 wags = 1.43643355948665e-07 pags = -7.15390916436254e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0530690668443025+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -6.47914036150301e-09 wvoff = -5.87717953730138e-08 pvoff = 1.92783322720727e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '6.94754145263125+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.89147912051856e-06 wnfactor = -7.97438389391246e-06 pnfactor = 3.35046114847282e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0247560778665857 leta0 = -2.1317982705245e-08 weta0 = -6.79850343887519e-08 peta0 = 6.09069236846211e-14
+ etab = 0.0105406711525826 letab = -5.3678367844527e-09 wetab = -3.69758449850672e-08 petab = 1.88299490586455e-14
+ dsub = 0.300865814793376 ldsub = -1.17608189390116e-08 wdsub = -7.74608790631168e-08 pdsub = 3.49748208919987e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.662413845611478 lpclm = 9.38158187847344e-08 wpclm = 9.21756931953574e-07 ppclm = -2.7913127515415e-13
+ pdiblc1 = 0.320534222962811 lpdiblc1 = 9.87277565172351e-08 wpdiblc1 = 4.05919528632457e-07 ppdiblc1 = -2.93759108218181e-13
+ pdiblc2 = 0.0192563236005596 lpdiblc2 = -2.21055121255114e-09 wpdiblc2 = -2.33435569089946e-08 ppdiblc2 = 6.57737576318046e-15
+ pdiblcb = -0.025
+ drout = 0.560273750149023 ldrout = -1.70865676908147e-07 wdrout = -3.82280541809809e-07 pdrout = 5.08401594893639e-13
+ pscbe1 = 354433812.358504 lpscbe1 = 54.0005132074944 wpscbe1 = 135.57973075314 ppscbe1 = -0.000160675611021187
+ pscbe2 = 1.6355008599768e-08 lpscbe2 = -2.00891715382625e-15 wpscbe2 = -8.48416768085536e-15 ppscbe2 = 5.9774245096837e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.74024680986435e-06 lalpha0 = 4.97466495995917e-12 walpha0 = 6.54015462506897e-11 palpha0 = -1.48018469564507e-17
+ alpha1 = 0.0
+ beta0 = 45.1022501519365 lbeta0 = -1.29225651086492e-06 wbeta0 = 7.27436586001246e-07 pbeta0 = 3.84503946622694e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.22443754820499e-08 lagidl = -4.20541580164323e-14 wagidl = -1.72472820812996e-13 pagidl = 1.1316214915752e-19
+ bgidl = 1225098106.98367 lbgidl = 425.972561563068 wbgidl = 1732.31029376787 pbgidl = -0.00126745835441258
+ cgidl = 1671.92003742666 lcgidl = -0.000810022886041529 wcgidl = -0.00342747586768102 pcgidl = 2.41017935618072e-9
+ egidl = 3.42724495190953 legidl = -1.86710646493062e-06 wegidl = -8.7662827549408e-06 pegidl = 5.55547446265195e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.815369136079391 lkt1 = -3.8108967740505e-07 wkt1 = -2.42234829815111e-06 pkt1 = 7.34074034831492e-13
+ kt2 = -0.019032
+ at = 40228.1945783334 lat = -0.00731239675301626 wat = 0.00772293499717636 pat = -1.58564431327679e-8
+ ute = -1.2463100961815 lute = -1.65602714283272e-07 wute = -8.65201761350892e-07 pute = 6.1364434923812e-13
+ ua1 = 5.534185e-10 lua1 = -7.2237112499977e-19
+ ub1 = -7.53108446284004e-19 lub1 = -2.01270365947307e-24 wub1 = -1.06536816367548e-23 pub1 = 7.55612370086835e-30
+ uc1 = -4.5116068918284e-10 luc1 = 2.42535618802929e-16 wuc1 = 5.04544531012064e-16 puc1 = -3.57848208620307e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.55 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1.5e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.479718076010656+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.24444837867179e-07 wvth0 = -3.16936381945268e-07 pvth0 = 1.80872481294687e-13
+ k1 = 0.439823410429467 lk1 = 4.39593526934539e-08 wk1 = 4.98591512721738e-07 pk1 = -1.77865361162549e-13
+ k2 = 0.102242166050673 lk2 = -2.36155421933232e-08 wk2 = -2.192180104795e-07 pk2 = 8.78656165066377e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -297531.869596497 lvsat = 0.190105268018834 wvsat = 0.497833957552635 pvsat = -2.56696435961201e-7
+ ua = 3.71254445317336e-09 lua = -1.23827388590308e-16 wua = -7.23101414376659e-15 pua = 1.97796407007115e-21
+ ub = -8.42707050214492e-18 lub = 3.52359078971755e-24 wub = 1.68879544396448e-23 pub = -6.83140838618726e-30
+ uc = 2.66361792467217e-10 luc = -1.36756113068655e-16 wuc = -3.9153560356749e-16 puc = 1.98960035015877e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00574979775194839 lu0 = 7.38806197388808e-09 wu0 = 5.9789996192277e-09 pu0 = -7.14858941432348e-15
+ a0 = 0.070361740752297 la0 = 3.94477121897393e-07 wa0 = 1.29890159628679e-06 pa0 = -6.63701301375068e-13
+ keta = -0.363101170008507 lketa = 1.67236020400735e-07 wketa = 4.39425361536022e-07 pketa = -2.36385016868278e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 5.53133506073384 lags = -2.4501435476961e-06 wags = -7.84508014716465e-06 pags = 3.99671835231683e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '0.27346164211768+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.72764903900393e-07 wvoff = -4.50819004303309e-07 pvoff = 2.18928373419826e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '6.54190656025194+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.6849095515744e-06 wnfactor = -3.27064255729318e-06 pnfactor = 9.55080872799448e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.01580269862506 leta0 = 5.08586574223126e-07 weta0 = 1.27507747659074e-06 peta0 = -6.23047660031683e-13
+ etab = 0.0664306462193101 letab = -3.38298065871837e-08 wetab = -1.36904918681211e-08 petab = 6.97188298384067e-15
+ dsub = 0.136256671460085 ldsub = 7.20663873034672e-08 wdsub = 1.89083057851627e-07 pdsub = -1.00762678981835e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.56090542718983 lpclm = -1.38224101913404e-06 wpclm = -3.23940473908767e-06 ppclm = 1.8399403058236e-12
+ pdiblc1 = 1.83533027189823 lpdiblc1 = -6.72682131403126e-07 wpdiblc1 = -8.42404808765055e-07 ppdiblc1 = 3.41950060601502e-13
+ pdiblc2 = 0.0605090135217994 lpdiblc2 = -2.32184835549425e-08 wpdiblc2 = -5.37577509649013e-08 ppdiblc2 = 2.2065804086151e-14
+ pdiblcb = 1.59860170066667 lpdiblcb = -8.26819166064502e-07 wpdiblcb = -2.39553663484184e-06 ppdiblcb = 1.21992703129321e-12
+ drout = -2.94796269644758 ldrout = 1.61570373352117e-06 wdrout = 3.13725228976994e-06 pdrout = -1.28392049958835e-12
+ pscbe1 = 727753101.983397 lpscbe1 = -136.112335033983 wpscbe1 = -589.767557204716 ppscbe1 = 0.000208707495371353
+ pscbe2 = 4.51575515409641e-09 lpscbe2 = 4.020222663382e-15 wpscbe2 = 1.40845215578492e-14 ppscbe2 = -5.5156804851266e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.88284439070776e-05 lalpha0 = -4.77676907876436e-11 walpha0 = -3.28289358041667e-11 palpha0 = 3.52220260299849e-17
+ alpha1 = -8.11800850333335e-10 lalpha1 = 4.13409583032251e-16 walpha1 = 1.19776831742092e-15 palpha1 = -6.09963515646603e-22
+ beta0 = 377.433352107628 lbeta0 = -0.000170531870181801 wbeta0 = -0.000472449140061111 pbeta0 = 2.44810211123769e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.50632919648105e-07 lagidl = 7.14461045285991e-14 wagidl = 3.52427484006659e-13 pagidl = -1.54143331071889e-19
+ bgidl = 7385190946.50168 lbgidl = -2711.05471696148 wbgidl = -9446.37141546862 pbgidl = 0.0044252853060161
+ cgidl = -3811.26191228474 lcgidl = 0.00198228752184901 wcgidl = 0.00986242242326289 pcgidl = -4.35770134848246e-9
+ egidl = -14.8688587072428 legidl = 7.45018432349273e-06 wegidl = 2.7176353502586e-05 pegidl = -1.27483130514936e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 1.7569876044078 lkt1 = -8.60608882401292e-07 wkt1 = -2.68635795050761e-06 pkt1 = 8.6852095029404e-13
+ kt2 = -0.019032
+ at = 5741.50281666659 lat = 0.0102499510266125 wat = 0.0364744964101606 pat = -3.04981757823301e-8
+ ute = -2.90505813892767 lute = 6.79114726485216e-07 wute = 2.05619650504028e-06 pute = -8.74077717921583e-13
+ ua1 = 5.52e-10
+ ub1 = -9.16382311598535e-18 lub1 = 2.27045278607234e-24 wub1 = 1.25157438236401e-23 pub1 = -4.24290621483777e-30
+ uc1 = 2.5099730656e-11 wuc1 = -1.98152000397473e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.56 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.946266572404+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = 4.16998994031929e-8
+ k1 = 0.57463991368 wk1 = 9.95938786049872e-9
+ k2 = 0.02677868733568 wk2 = -1.5112939312937e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 375817.673048 wvsat = -0.28840199632798
+ ua = 3.51442702460324e-09 wua = -1.23291312284281e-15
+ ub = -1.059473464076e-18 wub = 1.27501177195708e-24
+ uc = 1.8222228631144e-11 wuc = -6.17757859069069e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02153075062268 wu0 = -2.85624305783072e-9
+ a0 = 1.0637165987314 wa0 = -1.5342911941005e-7
+ keta = -0.0124276434096 wketa = 4.14149342592068e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.17092428540856 wags = -3.25095720191583e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.082107614352132+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' wvoff = -2.49446080986503e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.51932430484+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = 8.13820153121043e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.32078245010308 wpclm = -2.18231773413575e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -0.0029006459454072 wpdiblc2 = 6.18307179756727e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 205823461.64888 wpscbe1 = 18.4302214325066
+ pscbe2 = 1.495870890448e-08 wpscbe2 = 3.90315894186015e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.5867466425788e-05 walpha0 = 1.26915383848055e-10
+ alpha1 = 0.0
+ beta0 = 34.405916560192 wbeta0 = 4.51978897221495e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.13763790464e-08 wagidl = 2.23919277584947e-14
+ bgidl = 2323927891.6 wbgidl = -783.798067749654
+ cgidl = -1350.231344 wcgidl = 0.00268270216357943
+ egidl = -0.33330798459196 wegidl = 1.80773865143749e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.64463138316 wkt1 = -2.97256064842111e-7
+ kt2 = -0.019032
+ at = 713175.90816 wat = -0.54828445077104
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -5.0741587948e-18 wub1 = 1.94841319155248e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.57 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.946266572404+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = 4.16998994031925e-8
+ k1 = 0.57463991368 wk1 = 9.95938786049872e-9
+ k2 = 0.02677868733568 wk2 = -1.51129393129372e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 375817.673048 wvsat = -0.28840199632798
+ ua = 3.51442702460324e-09 wua = -1.23291312284281e-15
+ ub = -1.059473464076e-18 wub = 1.27501177195708e-24
+ uc = 1.8222228631144e-11 wuc = -6.17757859069069e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.02153075062268 wu0 = -2.85624305783072e-9
+ a0 = 1.0637165987314 wa0 = -1.53429119410049e-7
+ keta = -0.0124276434096 wketa = 4.14149342592068e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.17092428540856 wags = -3.25095720191583e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.082107614352132+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' wvoff = -2.49446080986503e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.51932430484+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = 8.13820153121045e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.32078245010308 wpclm = -2.18231773413575e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -0.0029006459454072 wpdiblc2 = 6.18307179756727e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 205823461.64888 wpscbe1 = 18.4302214325066
+ pscbe2 = 1.495870890448e-08 wpscbe2 = 3.90315894185889e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.5867466425788e-05 walpha0 = 1.26915383848055e-10
+ alpha1 = 0.0
+ beta0 = 34.405916560192 wbeta0 = 4.51978897221495e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.13763790464e-08 wagidl = 2.23919277584947e-14
+ bgidl = 2323927891.6 wbgidl = -783.798067749653
+ cgidl = -1350.231344 wcgidl = 0.00268270216357943
+ egidl = -0.33330798459196 wegidl = 1.80773865143749e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.644631383159999 wkt1 = -2.9725606484211e-7
+ kt2 = -0.019032
+ at = 713175.90816 wat = -0.54828445077104
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -5.0741587948e-18 wub1 = 1.94841319155248e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.58 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.970786039498579+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.93930595117797e-07 wvth0 = 7.78770490500205e-08 pvth0 = -2.86134120844174e-13
+ k1 = 0.613249194219438 lk1 = -3.05370452106546e-07 wk1 = -4.70065206742921e-08 pk1 = 4.50557612078795e-13
+ k2 = 0.0146578823728739 lk2 = 9.58664766520743e-08 wk2 = 1.63722992678587e-08 pk2 = -1.41445809510396e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 452224.009262194 lvsat = -0.60431681470211 wvsat = -0.401135419469867 pvsat = 8.9163682698497e-7
+ ua = 2.97337168670849e-09 lua = 4.27934193124408e-15 wua = -4.34615188767346e-16 pua = -6.31393793508637e-21
+ ub = -8.09805836481051e-19 lub = -1.97468368355535e-24 wub = 9.06640669492621e-25 pub = 2.91353914216701e-30
+ uc = 4.72154531599621e-11 luc = -2.29314661104555e-16 wuc = -1.04553723065053e-16 puc = 3.38341399468071e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0200931126121938 lu0 = 1.13706384344384e-08 wu0 = -7.35085805810822e-10 pu0 = -1.67767629955384e-14
+ a0 = 0.989509847529271 la0 = 5.86919746945435e-07 wa0 = -4.39410651758736e-08 pa0 = -8.65968392951654e-13
+ keta = -0.0155646236205401 lketa = 2.48111607333778e-08 wketa = 8.76993833023137e-09 pketa = -3.66075278594193e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.17158990940506 lags = -5.26458659431712e-09 wags = -3.34916642822981e-08 pags = 7.76761323223853e-15
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0618789272081338+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.59993743793667e-07 wvoff = -5.47909436305138e-08 pvoff = 2.36062129305392e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '1.06048455610196+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 1.15383282827063e-05 wnfactor = 2.96625942503758e-06 pnfactor = -1.70241803114059e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.453315568875e-05 lcit = -7.5400111631246e-11 wcit = -1.40656564283434e-11 pcit = 1.11248793105875e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.90346002666485 lpclm = -1.25177926224212e-05 wpclm = -4.51747303376351e-06 ppclm = 1.84693270535809e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00699621661092798 lpdiblc2 = 3.23928922862702e-08 wpdiblc2 = 1.22258651537272e-08 ppdiblc2 = -4.77939633522082e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 206473737.264721 lpscbe1 = -5.14319241458998 wpscbe1 = 17.4707748762166 ppscbe1 = 7.5885026753382e-6
+ pscbe2 = 1.49752317699197e-08 lpscbe2 = -1.30683473479319e-16 wpscbe2 = 1.46529936969822e-17 ppscbe2 = 1.92816408211155e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000188354295464569 lalpha0 = 9.68778952574979e-10 walpha0 = 3.07638085806009e-10 palpha0 = -1.42938103046094e-15
+ alpha1 = 1.90663113775e-10 lalpha1 = -1.50800223262492e-15 walpha1 = -2.81313128566869e-16 palpha1 = 2.22497586211751e-21
+ beta0 = -34.3080743828642 lbeta0 = 0.000543476132866367 wbeta0 = 0.000105903572053183 pbeta0 = -8.0186968633315e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.22607144789995e-09 lagidl = -9.9675931572042e-14 wagidl = 3.7976925864818e-15 pagidl = 1.47066454534243e-19
+ bgidl = 2232218933.87423 lbgidl = 725.34907389259 wbgidl = -648.48645290899 pbgidl = -0.00107021338967852
+ cgidl = -3081.452417077 lcgidl = 0.0136926602722343 wcgidl = 0.00523702537096659 pcgidl = -2.0202780828027e-8
+ egidl = 0.581998511225766 legidl = -7.23938790204636e-06 wegidl = 4.57253343409207e-07 pegidl = 1.06813259225227e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.502339501349717 lkt1 = -1.12542206620798e-06 wkt1 = -5.07200052691566e-07 pkt1 = 1.6604994858983e-12
+ kt2 = -0.019032
+ at = 843894.53896414 lat = -1.03388633068765 wat = -0.741152731716485 pat = 1.52544345106776e-6
+ ute = -1.27830384322982 lute = -2.19715925293451e-06 wute = -4.09873228321928e-07 pute = 3.24178983110521e-12
+ ua1 = 2.2096e-11
+ ub1 = -3.78356017765702e-18 lub1 = -1.02076671126381e-23 wub1 = 4.42046242833467e-26 pub1 = 1.50608616106734e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.59 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.864846289978916+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.20214370691941e-07 wvth0 = -7.54467241253751e-08 pvth0 = 3.13246839441738e-13
+ k1 = 0.51349360807869 lk1 = 8.45990730141704e-08 wk1 = 1.00177459874729e-07 pk1 = -1.24821363882466e-13
+ k2 = 0.0561869388909532 lk2 = -6.64809875412275e-08 wk2 = -4.19016219368717e-08 pk2 = 8.6361516959196e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 112957.541040318 lvsat = 0.721960626194257 wvsat = 0.0994339340022268 pvsat = -1.06521391807581e-6
+ ua = 3.48178012635833e-09 lua = 2.29184623854293e-15 wua = -1.18428917506341e-15 pua = -3.38327490415848e-21
+ ub = -1.16878759458449e-18 lub = -5.71334245689483e-25 wub = 1.32214013501967e-24 pub = 1.28924785655539e-30
+ uc = 5.77342299868566e-11 luc = -2.70435189415092e-16 wuc = -1.01858918807805e-16 puc = 3.27806735925421e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0208987552637788 lu0 = 8.22117989872948e-09 wu0 = -2.13078901631789e-09 pu0 = -1.13206102198636e-14
+ a0 = 1.56869513386951 la0 = -1.67726033368014e-06 wa0 = -7.57598195423818e-07 pa0 = 1.92389574347012e-12
+ keta = -0.204865052880046 lketa = 7.64833863816103e-07 wketa = 2.88072499479453e-07 pketa = -1.12847106503201e-12
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.21059565856311 lags = -4.06699781149045e-06 wags = -1.56788754944372e-06 pags = 6.00610472729952e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0824821094867173+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -7.94507534711149e-08 wvoff = -2.43920607503068e-08 pvoff = 1.17225296405942e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.2114938173305+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -4.68900467175136e-06 wnfactor = -2.87381406257952e-06 pnfactor = 5.80612697006128e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.04421768137306e-05 lcit = 2.22347069540764e-11 wcit = 2.27840980111116e-11 pcit = -3.28061094365643e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.0689896220399999 leta0 = 5.8243767995987e-07 weta0 = 2.1982614188043e-07 peta0 = -8.5935534514607e-13
+ etab = 0.0591591033464759 letab = -5.04915224757211e-07 wetab = -1.90567282396145e-07 petab = 7.44975148707128e-13
+ dsub = 0.00128891735000058 ldsub = 2.18414129984951e-06 wdsub = 8.24348032051612e-07 pdsub = -3.22258254429777e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.54494780980401 lpclm = -7.20702873865796e-06 wpclm = -2.51306161744505e-06 ppclm = 1.06335817243379e-11
+ pdiblc1 = 0.391691590921237 lpdiblc1 = -6.61285180884383e-09 wpdiblc1 = -2.49585105837482e-09 ppdiblc1 = 9.75690574995173e-15
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.705265198091947 ldrout = -5.67877975640943e-07 wdrout = -2.1433095546397e-07 pdrout = 8.37873287647526e-13
+ pscbe1 = 363168680.227529 lpscbe1 = -617.70289819195 wpscbe1 = -213.724151938488 ppscbe1 = 0.00091138727032572
+ pscbe2 = 1.44958057655718e-08 lpscbe2 = 1.74351263401788e-15 wpscbe2 = 7.22020174108138e-16 ppscbe2 = -2.57245874181115e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000654987888843972 lalpha0 = -2.32805648143319e-09 walpha0 = -9.36667766663291e-10 palpha0 = 3.43492162330467e-15
+ alpha1 = -3.8132622755e-10 lalpha1 = 7.28047099949837e-16 walpha1 = 5.62626257133737e-16 palpha1 = -1.07419418143259e-21
+ beta0 = 202.198098885013 lbeta0 = -0.000381085624981083 wbeta0 = -0.000243048515270213 pbeta0 = 5.62271261035839e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.29299212694755e-08 lagidl = 3.38483829583581e-14 wagidl = 4.80153447781911e-14 pagidl = -2.57914022961965e-20
+ bgidl = 3206601147.8926 lbgidl = -3083.75459625875 wbgidl = -1815.84409636932 pbgidl = 0.00349327947801878
+ cgidl = -992.757093792 lcgidl = 0.00552742807968238 wcgidl = 0.00112424794017403 pcgidl = -4.12490565670114e-9
+ egidl = -2.28099851112266 legidl = 3.95278320756925e-06 wegidl = 4.68145084804511e-06 pegidl = -5.83211817247522e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.618142983696716 lkt1 = -6.72717302842975e-07 wkt1 = -3.79396040662634e-07 pkt1 = 1.1608816518742e-12
+ kt2 = -0.019032
+ at = 342754.941029028 lat = 0.925193642540192 wat = 0.0687751602206268 pat = -1.64076716048739e-6
+ ute = -2.24017972938735 lute = 1.5630540550268e-06 wute = 8.03259496002821e-07 pute = -1.50064927146132e-12
+ ua1 = -7.26361199255202e-11 lua1 = 3.70331539818839e-16 wua1 = -6.07159803873747e-16 pua1 = 2.37353946329345e-21
+ ub1 = -5.7351885660459e-18 lub1 = -2.57826383532887e-24 wub1 = 3.62698979394673e-24 pub1 = 1.0548586861668e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.60 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.925075039512509+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.0522263064493e-07 wvth0 = 3.0647814425143e-08 pvth0 = 1.10685841714162e-13
+ k1 = 0.56275275317729 lk1 = -9.44894976533098e-09 wk1 = 2.74982512755803e-08 pk1 = 1.39414151354583e-14
+ k2 = 0.018509749003067 lk2 = 5.45418725221937e-09 wk2 = 6.0305628651484e-09 pk2 = -5.1530068740608e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 615647.688167738 lvsat = -0.23780053720877 wvsat = -0.602011754551337 pvsat = 2.74021262795079e-7
+ ua = 3.41067015273188e-09 lua = 2.42761295568923e-15 wua = -1.08099649533305e-15 pua = -3.58048645293367e-21
+ ub = -3.71121533524489e-19 lub = -2.09427817276829e-24 wub = 3.48530814671479e-25 pub = 3.14811145143018e-30
+ uc = -1.60221542248213e-10 luc = 1.45696868724714e-16 wuc = 1.35318318341354e-16 puc = -1.25023904101609e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0221967396338391 lu0 = 5.74300324019189e-09 wu0 = -3.41222135160667e-09 pu0 = -8.8740355337135e-15
+ a0 = 0.564678600023194 la0 = 2.3965823356594e-07 wa0 = 4.37362208328509e-07 pa0 = -3.57582407394005e-13
+ keta = 0.244413873626346 lketa = -9.29519266162268e-08 wketa = -3.74814295518698e-07 pketa = 1.37145548318205e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.872983012763503 lags = -8.89252332601019e-08 wags = 1.52691043448288e-06 pags = 9.73616764876726e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.112542685953607+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -2.20575978517055e-08 wvoff = 1.99606965554598e-08 pvoff = 3.25447945199075e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.33458194383074+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -3.01476067727194e-06 wnfactor = -1.02029926165833e-06 pnfactor = 2.26730383640248e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.24826912753876e-06 lcit = 6.59048870421462e-12 wcit = 1.06944296911506e-11 pcit = -9.72391019667864e-18
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.306212879403642 leta0 = -1.33917695921404e-07 weta0 = -3.33764888064586e-07 peta0 = 1.97588328776451e-13
+ etab = -0.205543336899806 letab = 4.67909283002908e-10 wetab = 1.99986874255471e-07 petab = -6.90374879969534e-16
+ dsub = 1.23025905219471 ldsub = -1.62269930102746e-07 wdsub = -9.88931037524474e-07 pdsub = 2.39420519290377e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.3572837250317 lpclm = 2.15255681922712e-06 wpclm = 4.71991929677254e-06 ppclm = -3.17598708613199e-12
+ pdiblc1 = 0.271758261939298 lpdiblc1 = 2.22369856549922e-07 wpdiblc1 = 1.7445929945471e-07 ppdiblc1 = -3.28094715367156e-13
+ pdiblc2 = 0.00257196283119567 lpdiblc2 = -2.44758753546034e-09 wpdiblc2 = -1.89146693143633e-09 ppdiblc2 = 3.61128323884481e-15
+ pdiblcb = -0.025
+ drout = 1.04996238088609 ldrout = -1.22599107189065e-06 wdrout = -7.22913035028851e-07 pdrout = 1.80888362305677e-12
+ pscbe1 = 41649287.2565508 lpscbe1 = -3.84199716210901 wpscbe1 = 260.660350342971 ppscbe1 = 5.66865934484534e-6
+ pscbe2 = 1.47890132863298e-08 lpscbe2 = 1.18370617501071e-15 wpscbe2 = 2.8940831043586e-16 ppscbe2 = -1.74649454109486e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000999909737729803 lalpha0 = 8.31556812102793e-10 walpha0 = 1.50504431687448e-09 palpha0 = -1.22691717218982e-15
+ alpha1 = 0.0
+ beta0 = -6.96579482348511 lbeta0 = 1.82605390818674e-05 wbeta0 = 6.55615150464158e-05 pbeta0 = -2.69424393461849e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.4296307767941e-08 lagidl = 3.64571563805534e-14 wagidl = 7.0862460098252e-14 pagidl = -6.94122572210228e-20
+ bgidl = 1527883643.4601 lbgidl = 121.336799079005 wbgidl = 131.329568767718 pbgidl = -0.000224361842144116
+ cgidl = 2725.44660408318 lcgidl = -0.00157155233048581 wcgidl = -0.00141358734229611 pcgidl = 7.20456356354983e-10
+ egidl = -2.61790291183535 legidl = 4.59601793462995e-06 wegidl = 5.17853509845904e-06 pegidl = -6.78117627757802e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.749671378285862 lkt1 = -4.21596715473647e-07 wkt1 = -7.93014036239782e-08 pkt1 = 5.87925966108143e-13
+ kt2 = -0.019032
+ at = 1605982.98471986 lat = -1.48662449987654 wat = -1.56180254081974 pat = 1.47241331522392e-6
+ ute = -1.554081257815 lute = 2.53120548177288e-07 wute = 1.87389768483609e-07 pute = -3.24799994195269e-13
+ ua1 = -2.70618672148961e-10 lua1 = 7.48329727651442e-16 wua1 = 1.2143196077475e-15 pua1 = -1.10412010334441e-21
+ ub1 = -1.0263146780052e-17 lub1 = 6.06674038476229e-24 wub1 = 7.97968895025961e-24 pub1 = -7.25553217802355e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.61 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.52463471660839+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 4.39927005754504e-07 wvth0 = 6.92761834901119e-07 pvth0 = -4.9134133140362e-13
+ k1 = 0.465125555305598 lk1 = 7.93185798995032e-08 wk1 = 1.94721000538898e-07 pk1 = -1.38105869632214e-13
+ k2 = -0.00487320855871004 lk2 = 2.67151414152651e-08 wk2 = 1.65141205537685e-09 pk2 = -1.17126400027602e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1408317.12091373 lvsat = -0.958535218933063 wvsat = -1.36678962515362 pvsat = 9.69395541640203e-7
+ ua = 2.27437497585534e-08 lua = -1.5150989675904e-14 wua = -2.28169125815762e-14 pua = 1.61828952484829e-20
+ ub = -1.50983015356272e-17 lub = 1.12964102441436e-23 wub = 1.73250654733511e-23 pub = -1.22878026869743e-29
+ uc = 6.77923030150765e-12 luc = -6.1485837161193e-18 wuc = -9.92861574866739e-18 puc = 7.04187071974235e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0733522117613004 lu0 = -4.07701097917023e-08 wu0 = -5.98829889883094e-08 pu0 = 4.24720099399584e-14
+ a0 = 0.942610790685141 la0 = -1.03976610793438e-07 wa0 = 2.00445902643454e-07 pa0 = -1.42166256449869e-13
+ keta = 0.875554976142642 lketa = -6.66816974079169e-07 wketa = -1.01827174941085e-06 pketa = 7.22209238269648e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -7.02252933270158 lags = 5.5025497581436e-06 wags = 7.42852494520614e-06 pags = -5.26868131738746e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.325415190732614+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.71496727118606e-07 wvoff = 2.53470289314796e-07 pvoff = -1.79773802696519e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '-2.73558008296921+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 3.41378414559591e-06 wnfactor = 6.69798366369825e-06 pnfactor = -4.75054491347799e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.273125e-05 lcit = 1.61221390625e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.69833150413179 leta0 = -4.90451555455472e-07 weta0 = -5.29436978481369e-07 peta0 = 3.75503176987911e-13
+ etab = -0.917591728340729 letab = 6.47897909200663e-07 wetab = 9.0573845268409e-07 petab = -6.42394997566191e-13
+ dsub = 3.84122942635146 ldsub = -2.53629474280477e-06 wdsub = -3.29882513289375e-06 pdsub = 2.3396917255049e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.04171203503977 lpclm = 3.68412326010196e-06 wpclm = 5.57799767229219e-06 ppclm = -3.95619484907323e-12
+ pdiblc1 = 0.736857725441143 lpdiblc1 = -2.00521830639131e-07 wpdiblc1 = -8.47337986689803e-07 ppdiblc1 = 6.00974467059743e-13
+ pdiblc2 = -0.0239630975856034 lpdiblc2 = 2.16794161485142e-08 wpdiblc2 = 9.45733465718165e-09 ppdiblc2 = -6.70761460560609e-15
+ pdiblcb = -0.025
+ drout = -3.29316526542489 ldrout = 2.7229977405176e-06 wdrout = 5.75787472978396e-06 pdrout = -4.08377265209927e-12
+ pscbe1 = -1138144250.84545 lpscbe1 = 1068.88527735714 wpscbe1 = 1213.37041447096 ppscbe1 = -0.000860582966463527
+ pscbe2 = 2.53341744242803e-08 lpscbe2 = -8.40448158967084e-15 wpscbe2 = -7.41675017415522e-15 ppscbe2 = 5.2603300610196e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000503151529201403 lalpha0 = 3.79879410998345e-10 walpha0 = 7.07721864641514e-10 palpha0 = -5.01951732496994e-16
+ alpha1 = 0.0
+ beta0 = -108.626614991932 lbeta0 = 0.000110695639820028 wbeta0 = 0.000163346841048844 pbeta0 = -1.15853747013892e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.1496057212765e-08 lagidl = -5.17955147815358e-15 wagidl = -2.49028268834358e-14 pagidl = 1.76623299670768e-20
+ bgidl = 1210002259.4755 lbgidl = 410.370447467001 wbgidl = -524.752158710337 pbgidl = 0.000372180468565308
+ cgidl = 2724.2124713841 lcgidl = -0.00157043019532917 wcgidl = -0.00282423967313879 pcgidl = 2.00309198817368e-9
+ egidl = 10.5035421773808 legidl = -7.33465601273982e-06 wegidl = -1.03629661965207e-05 pegidl = 7.3499337748823e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -3.16772621215034 lkt1 = 1.77701964221763e-06 wkt1 = 2.57910582431521e-06 pkt1 = -1.82923080589556e-12
+ kt2 = -0.019032
+ at = -202847.3551 lat = 0.158054486604675 wat = 0.261721774917875 pat = -1.85626168860503e-7
+ ute = -0.551898427455004 lute = -6.58114190327542e-07 wute = -7.72079236007731e-07 pute = 5.47597198138482e-13
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.62 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.9293834525+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.7745046685624e-8
+ k1 = 0.4486544625 lk1 = 9.10007024718747e-8
+ k2 = 0.0545935165462499 lk2 = -1.54616333654278e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 19390.418875 lvsat = 0.0265610444879062
+ ua = 1.84212674625e-09 lua = -3.26513554427813e-16
+ ub = 7.85113574999999e-19 lub = 3.10980769312502e-26
+ uc = 3.10172318250001e-13 luc = -1.56040434149381e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.01860092625 lu0 = -1.93776054281249e-9
+ a0 = 0.678882499999999 la0 = 8.30726793750007e-8
+ keta = -0.0980569012499999 lketa = 2.37172499615625e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.770199644674999 lags = -2.44432690607436e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0929023073512499+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 6.58696458037406e-9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '1.54281373375+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 3.79333331087812e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.02132153825 leta0 = 1.99623648538125e-8
+ etab = -0.014520120625 letab = 7.39437142828125e-9
+ dsub = 0.24836583915 ldsub = 1.19437564178627e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.28714489775 lpclm = -9.53685194791875e-8
+ pdiblc1 = 0.595650715625 lpdiblc1 = -1.00370758927032e-7
+ pdiblc2 = 0.00343496727237499 lpdiblc2 = 2.24733864799303e-9
+ pdiblcb = -0.025
+ drout = 0.3011788447375 ldrout = 1.73709180384928e-7
+ pscbe1 = 446324488.6375 lpscbe1 = -54.8991761211469
+ pscbe2 = 1.06047692275e-08 lpscbe2 = 2.04234904614563e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.958638137625e-05 lalpha0 = -5.05745207885529e-12
+ alpha1 = 0.0
+ beta0 = 45.59527842 lbeta0 = 1.31376191761501e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -4.46510045e-08 lagidl = 3.4642752041625e-14 wagidl = 1.26217744835362e-29 pagidl = 6.01853107621011e-36
+ bgidl = 2399190750 lbgidl = -433.061489437501
+ cgidl = -651.090000000001 lcgidl = 0.0008235030825
+ egidl = -2.5142010616625 legidl = 1.89817837955163e-06 wegidl = -2.11758236813575e-22 pegidl = -4.03896783473158e-28
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.826404468749998 lkt1 = 1.16437195710938e-7
+ kt2 = -0.019032
+ at = 45462.5 lat = -0.018059278125
+ ute = -1.83271025 lute = 2.503015948125e-7
+ ua1 = 5.53418499999999e-10 lua1 = -7.22371125000165e-19
+ ub1 = -7.97376012499999e-18 lub1 = 3.10854354365625e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.63 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 1e-06 wmax = 1.5e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.731347573152121+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -8.3104724872282e-08 wvth0 = 5.43293530941169e-08 pvth0 = -2.76672230631788e-14
+ k1 = 0.529206660873701 lk1 = 4.99794954500678e-08 wk1 = 3.66711353386794e-07 pk1 = -1.86747756712225e-13
+ k2 = -0.00411231214659974 lk2 = 1.4434309896406e-08 wk2 = -6.22977210412471e-08 pk2 = 3.17251144402551e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 324236.512453956 lvsat = -0.128681828667177 wvsat = -0.419551714670178 pvsat = 2.13656710695788e-7
+ ua = -5.19344031931497e-09 lua = 3.25634897371115e-15 wua = 5.90928546486223e-15 pua = -3.00930362298109e-21
+ ub = 9.5181654609053e-18 lub = -4.41620859596602e-24 wub = -9.58927218109383e-24 pub = 4.88333685822203e-30
+ uc = -1.72065167409975e-11 luc = 7.35996956192797e-18 wuc = 2.68541239805337e-17 puc = -1.36754626370868e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00694536733226694 lu0 = 3.99783283604309e-09 wu0 = 4.21500126422512e-09 pu0 = -2.14648939380665e-15
+ a0 = 0.194539743947901 la0 = 3.29724227894531e-07 wa0 = 1.11568365818385e-06 pa0 = -5.68161902930124e-13
+ keta = 0.251095277846505 lketa = -1.54088497243332e-07 wketa = -4.66788330665864e-07 pketa = 2.37711957391591e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -5.61837645448228 lags = 3.2289391094351e-06 wags = 8.60571710911492e-06 pags = -4.38246143781678e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.203861609677007+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 6.30929892897659e-08 wvoff = 2.53445678264156e-07 pvoff = -1.29067211656021e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.91425506187281+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -3.19073165258725e-07 wnfactor = 2.08176133538432e-06 pnfactor = -1.06013696004447e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.992012755e-05 lcit = 2.03293249548375e-11 wcit = 5.88999925131373e-11 pcit = -2.99948211873152e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.623955551515889 leta0 = -3.08644993109466e-07 weta0 = -1.14429727454673e-06 peta0 = 5.82733387062922e-13
+ etab = 0.08125553551469 letab = -4.13793814608559e-08 wetab = -3.55638154794323e-08 petab = 1.81108730329009e-14
+ dsub = 0.300894506263302 ldsub = -1.48064673095866e-08 wdsub = -5.38311769574418e-08 pdsub = 2.74135268655772e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.78215644629306 lpclm = 1.46767318997474e-06 wpclm = 4.64399452989518e-06 ppclm = -2.36495421434912e-12
+ pdiblc1 = 0.831833650779935 lpdiblc1 = -2.20646918654682e-07 wpdiblc1 = 6.38200266877447e-07 ppdiblc1 = -3.2500348590734e-13
+ pdiblc2 = 0.00966171079169956 lpdiblc2 = -9.23630489222993e-10 wpdiblc2 = 2.12646984590136e-08 ppdiblc2 = -1.08290476902527e-14
+ pdiblcb = -1.621805102 lpdiblcb = 8.13172998193499e-07 wpdiblcb = 2.35599970052549e-06 ppdiblcb = -1.19979284749261e-12
+ drout = -0.821654929325002 ldrout = 7.45512279826257e-7
+ pscbe1 = 3992032757.91542 lpscbe1 = -1860.55111225093 wpscbe1 = -5406.035918431 ppscbe1 = 0.00275302379146099
+ pscbe2 = -5.830437739442e-08 lpscbe2 = 3.71343319633584e-14 wpscbe2 = 1.06772234846028e-13 ppscbe2 = -5.43737605953396e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.67097169415412e-05 lalpha0 = 3.37963359894799e-11 walpha0 = 1.67150301467285e-10 palpha0 = -8.51212910222148e-17
+ alpha1 = 0.0
+ beta0 = -5.64479187731126 lbeta0 = 2.74077677165207e-05 wbeta0 = 9.2761975168892e-05 pbeta0 = -4.72390358547583e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.52950686440029e-07 lagidl = -6.59859090695849e-14 wagidl = -9.54937332616542e-14 pagidl = 4.86301836634974e-20
+ bgidl = 3850669213.192 lbgidl = -1172.22689681802 wbgidl = -4231.37546214378 pbgidl = 0.00215482795409672
+ cgidl = 1276.299898 lcgidl = -0.000158020223056503 wcgidl = 0.00235599970052549 pcgidl = -1.19979284749261e-9
+ egidl = -0.497156799849904 legidl = 8.70998589223562e-07 wegidl = 5.97168341013074e-06 pegidl = -3.04107977660908e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.75666108322903 lkt1 = -6.89738936634383e-07 wkt1 = -1.21043018614048e-06 pkt1 = 6.1641157229204e-13
+ kt2 = -0.019032
+ at = -1473.60203999997 lat = 0.00584293183886997 wat = 0.0471199940105098 pat = -2.39958569498521e-8
+ ute = -0.882306789812006 lute = -2.33691367288239e-07 wute = -9.28263882007044e-07 pute = 4.72718381912087e-13
+ ua1 = 5.52e-10
+ ub1 = -6.81138000000002e-19 lub1 = -6.05224273500002e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.64 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.959843529224+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = 5.49434876254343e-8
+ k1 = 0.62498167272 wk1 = -3.9146279628033e-8
+ k2 = 0.016196245398984 wk2 = 8.81130672608864e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -210585.346096 wvsat = 0.283602483083959
+ ua = 2.00680665770416e-09 wua = 2.37689133567428e-16
+ ub = 6.90279836712e-19 wub = -4.31778086283373e-25
+ uc = -8.1292615534288e-11 wuc = 3.52955707748871e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.01695872034616 wu0 = 1.60352558727963e-9
+ a0 = 0.9927399307044 wa0 = -8.41952124897841e-8
+ keta = -0.0095869438128 wketa = 1.37054436702051e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.17588942434192 wags = -3.73527969311484e-8
+ b0 = -8.29213795839999e-09 wb0 = 8.08853280296944e-15
+ b1 = -9.57066398879999e-11 wb1 = 9.335665905219e-17
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.10375224615976+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' wvoff = -3.83143858042676e-9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.64277997352+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = 6.93395814929808e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -9.50891999999999e-06 wcit = 1.415266797832e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.56120909605 wpclm = 2.57980139159309e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0096712918908144 wpdiblc2 = -6.08017467702374e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 222156089.19184 wpscbe1 = 2.49862522623641
+ pscbe2 = 1.5011313840776e-08 wpscbe2 = -1.22816852715827e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000195588957154592 walpha0 = -1.28121238707732e-10
+ alpha1 = 0.0
+ beta0 = 42.965495993128 wbeta0 = -3.82961854732472e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.46024021816e-08 wagidl = 4.5047659121633e-14
+ bgidl = 993726204.0 wbgidl = 513.741847613015
+ cgidl = 1980.3568 wcgidl = -0.0005661067191328
+ egidl = 2.7701879881744 wegidl = -1.21955408121356e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.83471880732 wkt1 = 8.63609952705064e-7
+ kt2 = -0.019032
+ at = -430282.4244 wat = 0.567097405891282
+ ute = -1.9788899288 wute = 4.12408744888244e-7
+ ua1 = 2.2096e-11
+ ub1 = -5.0409175896e-18 wub1 = 1.91598819090496e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.65 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.996968579329411+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 7.39131903811137e-07 wvth0 = 9.11569692505559e-08 pvth0 = -7.20983259044964e-13
+ k1 = 0.651432625425055 lk1 = -5.26618630143116e-07 wk1 = -6.49477556403685e-08 pk1 = 5.13688036298582e-13
+ k2 = 0.0102424878594144 lk2 = 1.18534847294677e-07 wk2 = 1.46188757030317e-08 pk2 = -1.15624342654203e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -402214.178730148 lvsat = 3.81518633612142 wvsat = 0.470526061361608 pvsat = -3.7215082508243e-6
+ ua = 1.84620125432388e-09 lua = 3.19753312724885e-15 wua = 3.9435103187311e-16 pua = -3.11902089884239e-21
+ ub = 9.82030211150698e-19 lub = -5.80853114229366e-24 wub = -7.16364822028104e-25 pub = 5.66590846862578e-30
+ uc = -1.05141662803544e-10 luc = 4.74816644345427e-16 wuc = 5.85590285374933e-17 puc = -4.63157996460169e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0158752258257738 lu0 = 2.15715632799983e-08 wu0 = 2.66041598321223e-09 pu0 = -2.10418951152213e-14
+ a0 = 1.04963023049076 la0 = -1.13264320102151e-06 wa0 = -1.39688627855186e-07 pa0 = 1.10483227986363e-12
+ keta = -0.0105130140441657 lketa = 1.84373637538176e-08 wketa = 2.27387586992525e-09 pketa = -1.79846527242063e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.201128529422031 lags = -5.02491652816196e-07 wags = -6.19721810251222e-08 pags = 4.90153472772948e-13
+ b0 = -1.37575206373562e-08 lb0 = 1.0881167010101e-13 wb0 = 1.34197184756266e-14 pb0 = -1.0613990835335e-19
+ b1 = -1.58787285015847e-10 lb1 = 1.25588833401159e-15 wb1 = 1.54888422019568e-16 pb1 = -1.22505125185827e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.101163361554475+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.15427508277677e-08 wvoff = -6.35675571311343e-09 pvoff = 5.02771701239424e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.17425575919192+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 9.32796571411127e-06 wnfactor = 1.15041588569928e-06 pnfactor = -9.09892684396699e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.90718096258333e-05 lcit = 1.90389960283122e-10 wcit = 2.34807504122806e-11 pcit = -1.8571512519833e-16
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.30436847788299 lpclm = 3.47049959227585e-05 wpclm = 4.28015923796455e-06 ppclm = -3.38528494528711e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0137796366517622 lpdiblc2 = -8.17940629319002e-08 wpdiblc2 = -1.00876431407112e-08 ppdiblc2 = 7.97856915106703e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 220467780.154178 lpscbe1 = 33.6129667080641 wpscbe1 = 4.14547952378734 ppscbe1 = -3.27876339235155e-5
+ pscbe2 = 1.50196125163933e-08 lpscbe2 = -1.65220407533688e-16 wpscbe2 = -2.03765952077753e-17 ppscbe2 = 1.61163585647168e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000282159861408401 lalpha0 = -1.72356177551514e-09 walpha0 = -2.12566480978493e-10 palpha0 = 1.68124143967914e-15
+ alpha1 = 0.0
+ beta0 = 45.553150810807 lbeta0 = -5.15182666788749e-05 wbeta0 = -6.35373608861041e-06 pbeta0 = 5.02532871588419e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.50408886028349e-08 lagidl = 6.06007435781972e-13 wagidl = 7.47387589472809e-14 pagidl = -5.91127529203781e-19
+ bgidl = 646593310.582251 lbgidl = 6911.15555827733 wbgidl = 852.351239965786 pbgidl = -0.00674145904469938
+ cgidl = 2362.87238503333 lcgidl = -0.00761559841132489 wcgidl = -0.000939230016491224 pcgidl = 7.42860500793321e-9
+ egidl = 3.59423481024676 legidl = -1.64061541923442e-05 wegidl = -2.02336725761676e-06 pegidl = 1.60033174823054e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -2.41825589517797 lkt1 = 1.16177857664364e-05 wkt1 = 1.43281887090777e-06 pkt1 = -1.13325226547273e-11
+ kt2 = -0.019032
+ at = -813467.41170714 lat = 7.6289257085447 wat = 0.940873669020084 pat = -7.44160506669709e-6
+ ute = -2.25755253249678 lute = 5.54796344265017e-06 wute = 6.84229067013856e-07 pute = -5.41173874827934e-12
+ ua1 = 2.2096e-11
+ ub1 = -6.33554158714531e-18 lub1 = 2.5774992823129e-23 wub1 = 3.17882399081455e-24 pub1 = -2.51421136493499e-29
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.66 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.799429444718611+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -8.23254496609319e-07 wvth0 = -8.927205590172e-08 pvth0 = 7.06075008140678e-13
+ k1 = 0.468410253525961 lk1 = 9.20951064799799e-07 wk1 = 9.42760446693979e-08 pk1 = -7.45652806301435e-13
+ k2 = 0.0582991279433052 lk2 = -2.61557133288836e-07 wk2 = -2.61973791588362e-08 pk2 = 2.07201621112025e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 211488.47937806 lvsat = -1.03874141252092 wvsat = -0.166310909786508 pvsat = 1.31539456322894e-6
+ ua = 3.57073354363451e-09 lua = -1.04422238819813e-14 wua = -1.01730942265841e-15 pua = 8.04615455116106e-21
+ ub = -6.84306541793995e-19 lub = 7.37094282093416e-24 wub = 7.84222884487311e-25 pub = -6.20261484913126e-30
+ uc = -6.77319227841574e-11 luc = 1.78933658097097e-16 wuc = 7.57123501013417e-18 puc = -5.98827905039036e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.023084479928291 lu0 = -3.54482297303358e-08 wu0 = -3.65300308882863e-09 pu0 = 2.88925146803179e-14
+ a0 = 0.970482533749587 la0 = -5.06644280571427e-07 wa0 = -2.53809480587364e-08 pa0 = 2.0074426343356e-13
+ keta = -0.000534772696822755 lketa = -6.04830416226547e-08 wketa = -5.890869633905e-09 pketa = 4.65923606519631e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.0988408611085875 lags = 3.06527087791905e-07 wags = 3.74711038823028e-08 pags = -2.96368328381104e-13
+ b0 = 8.1040100784688e-09 lb0 = -6.40966417131294e-14 wb0 = -7.90502421500208e-15 pb0 = 6.25228127725052e-20
+ b1 = 9.3535295495541e-11 lb1 = -7.39794035898108e-16 wb1 = -9.12386298499435e-17 pb1 = 7.21629133140666e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.151976274263611+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 3.50349279016964e-07 wvoff = 3.30941531653632e-08 pvoff = -2.61749930923148e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '6.9660321139803+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -2.85713914199987e-05 wnfactor = -2.79428331810462e-06 pnfactor = 2.21006853337189e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.13437499999997e-07 lcit = 3.8649044453125e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.497086103674554 lpclm = 4.59224780455046e-06 wpclm = -2.24977913108458e-07 ppclm = 1.77940655925307e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0055373989390125 lpdiblc2 = -1.66041443023346e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225920465.073143 lpscbe1 = -9.51368148725487 wpscbe1 = -1.49845797759735 ppscbe1 = 1.18516787593129e-5
+ pscbe2 = 1.49533720830446e-08 lpscbe2 = 3.58691739929416e-16 wpscbe2 = 3.59759378205929e-17 ppscbe2 = -2.84542686207546e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000180849902470727 lalpha0 = -9.22275982787351e-10 walpha0 = -5.25006722531846e-11 palpha0 = 4.152409420185e-16
+ alpha1 = -3.8132622755e-10 lalpha1 = 3.01600446524984e-15 walpha1 = 2.76631586471237e-16 palpha1 = -2.18794837529763e-21
+ beta0 = 172.630513426203 lbeta0 = -0.0010566048969447 wbeta0 = -9.59538456708203e-05 pbeta0 = 7.58922953871935e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.1508156093505e-08 lagidl = -1.57623095982555e-13 wagidl = -2.57408457527351e-14 pagidl = 2.0359078426982e-19
+ bgidl = 2218542799.7048 lbgidl = -5521.78593856518 wbgidl = -635.146122537961 pbgidl = 0.00502352946968337
+ cgidl = 4295.252191054 lcgidl = -0.0228992733920939 wcgidl = -0.00195855163221636 pcgidl = 1.54906744971073e-8
+ egidl = -1.53256546967815 legidl = 2.41429909216519e-05 wegidl = 2.51989632032601e-06 pegidl = -1.99304899715385e-11
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.368691307366637 lkt1 = -4.59273294971042e-06 wkt1 = -6.37566648919584e-07 pkt1 = 5.04267401796722e-12
+ kt2 = -0.019032
+ at = 457835.275913145 lat = -2.42612507351604 wat = -0.364572767810444 pat = 2.88349716380475e-6
+ ute = -1.69849443125 lute = 1.12623315536406e-6
+ ua1 = 2.2096e-11
+ ub1 = -3.73824283125e-18 lub1 = 5.23230763806405e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.67 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.02007147576571+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 3.92903632615677e-08 wvth0 = 7.59670624496152e-08 pvth0 = 6.01139847257244e-14
+ k1 = 0.71630439206244 lk1 = -4.81290962739339e-08 wk1 = -9.76535081190842e-08 pk1 = 4.64779793693757e-15
+ k2 = -0.0128117804976345 lk2 = 1.64331855339072e-08 wk2 = 2.54029028958487e-08 pk2 = 5.48321848974813e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -78637.0076552859 lvsat = 0.0954316476641868 wvsat = 0.286324070149159 pvsat = -4.54068732084569e-7
+ ua = 1.23409434694359e-09 lua = -1.30771710231728e-15 wua = 1.00820692772358e-15 pua = 1.27904758430245e-22
+ ub = -5.19012452076701e-19 lub = 6.72476690070682e-24 wub = 6.88319571361017e-25 pub = -5.8277048222923e-30
+ uc = -4.79207386264372e-12 luc = -6.71139462993304e-17 wuc = -4.08678858230249e-17 puc = 1.29477842613124e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0113679083377098 lu0 = 1.0354777760144e-08 wu0 = 7.16603749432844e-09 pu0 = -1.3401819719389e-14
+ a0 = 0.165933125620294 la0 = 2.63854049315802e-06 wa0 = 6.10720394474845e-07 pa0 = -2.28593490986585e-12
+ keta = 0.293593566378887 lketa = -1.21030425115437e-06 wketa = -1.98146966842196e-07 pketa = 7.98169508663475e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.05579318418875 lags = 4.82028022937052e-06 wags = 6.42852381663216e-07 pags = -2.66295508854614e-12
+ b0 = 1.68583618134721e-07 lb0 = -6.91451549507035e-13 wb0 = -1.64444215975041e-13 pb0 = 6.74473648160439e-19
+ b1 = 8.93551485454018e-10 lb1 = -3.86725732649328e-15 wb1 = -8.7161122228018e-16 pb1 = 3.77230069009857e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0107594551459677+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -2.01702571118683e-07 wvoff = -9.43536370363738e-08 pvoff = 2.36475342922992e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '-1.93884314876307+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 6.23999220088081e-06 wnfactor = 4.10095352964858e-06 pnfactor = -4.85451931336029e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.13754336274612e-05 lcit = -4.44694139081529e-11 wcit = -8.25226282330725e-12 pcit = 3.22601584420139e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.32257693306 leta0 = -9.48293875564805e-07 weta0 = -1.62125888025645e-07 peta0 = 6.33790627764252e-13
+ etab = -0.134410118122952 letab = 2.5179525427215e-07 wetab = -1.75095959067695e-09 petab = 6.84493877985391e-15
+ dsub = 1.00139128243825 ldsub = -1.72550887087171e-06 wdsub = -1.51197819564257e-07 pdsub = 5.91070076131574e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.52252635445367 lpclm = 1.25102001049087e-05 wpclm = 2.42998578618345e-06 ppclm = -8.59951028220381e-12
+ pdiblc1 = 0.820471817134348 lpdiblc1 = -1.68282195113245e-06 wpdiblc1 = -4.20747807597049e-07 ppdiblc1 = 1.64480836684876e-12
+ pdiblc2 = 0.00334169882537969 lpdiblc2 = -8.02060363311553e-09 wpdiblc2 = -2.00132141242131e-09 ppdiblc2 = 7.82366573150801e-15
+ pdiblcb = -0.025
+ drout = -0.10216486022926 ldrout = 2.58856797985124e-06 wdrout = 5.73273465205218e-07 pdrout = -2.2410692938535e-12
+ pscbe1 = 52996996.6449871 lpscbe1 = 666.487387465514 wpscbe1 = 88.8315761253693 ppscbe1 = -0.000341271007057711
+ pscbe2 = 1.46063095159276e-08 lpscbe2 = 1.71544608043147e-15 wpscbe2 = 6.14229732838565e-16 ppscbe2 = -2.54508133438151e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.00129869453818571 lalpha0 = 4.86163312184881e-09 walpha0 = 9.69043942053101e-10 palpha0 = -3.57823234145835e-15
+ alpha1 = 1.0396640102e-09 lalpha1 = -2.53900162167435e-15 walpha1 = -8.23472986318549e-16 palpha1 = 2.11263542588084e-21
+ beta0 = -388.704512187547 lbeta0 = 0.00113779405193586 wbeta0 = 0.000333345073090071 pbeta0 = -9.19313844294081e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -9.20053009303781e-08 lagidl = 3.2522188588806e-13 wagidl = 1.056401875669e-13 pagidl = -3.10010520234963e-19
+ bgidl = -1555853333.8917 lbgidl = 9233.27214669693 wbgidl = 2829.67307806925 pbgidl = -0.00852131499029037
+ cgidl = -1556.718474778 lcgidl = -2.24570666901049e-05 wcgidl = 0.0016743618134113 pcgidl = 1.28870760978731e-9
+ egidl = 6.16859773506181 legidl = -5.96278133647779e-06 wegidl = -3.56067401191055e-06 pegidl = 3.83997959975729e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.78359382060063 lkt1 = 9.38474700149582e-07 wkt1 = 7.57438316391948e-07 pkt1 = -4.10749142676882e-13
+ kt2 = -0.019032
+ at = -284475.971318125 lat = 0.475755169722804 wat = 0.680605044746009 pat = -1.20236419993156e-6
+ ute = -1.544125840346 lute = 5.22767741372601e-07 wute = 1.24296514152994e-07 pute = -4.85906147952592e-13
+ ua1 = -1.30716412814896e-09 lua1 = 5.19641015596632e-15 wua1 = 5.97055603635775e-16 pua1 = -2.33403961851315e-21
+ ub1 = -4.20529119779e-18 lub1 = 7.05811646496056e-24 wub1 = 2.13465752567099e-24 pub1 = -8.34490993222931e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.68 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.02799464789783+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 5.44176796548074e-08 wvth0 = 1.3104033474617e-07 pvth0 = -4.50346604064755e-14
+ k1 = 0.68119793884542 lk1 = 1.8897899530662e-08 wk1 = -8.80386313036548e-08 pk1 = -1.37094056229206e-14
+ k2 = -0.00342421692820261 lk2 = -1.49002021103062e-09 wk2 = 2.74259621969416e-08 pk2 = 1.62069251913654e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -34113.59686402 lvsat = 0.0104253256109622 wvsat = 0.0317952918877518 pvsat = 3.1890337811023e-8
+ ua = 3.08901387003978e-09 lua = -4.84922220178869e-15 wua = -7.67238161006176e-16 pua = 3.51767329408753e-21
+ ub = 7.79453424105219e-19 lub = 4.24567092660649e-24 wub = -7.7379292544859e-25 pub = -3.03616653775855e-30
+ uc = -7.57602766297423e-11 luc = 6.83820948337526e-17 wuc = 5.2930914638879e-17 puc = -4.96075171687665e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0231230638400158 lu0 = -1.20887528826337e-08 wu0 = -4.31580059322486e-09 pu0 = 8.5198796492722e-15
+ a0 = 1.80729777746693 la0 = -4.95234968380179e-07 wa0 = -7.74745697832276e-07 pa0 = 3.59266226871527e-13
+ keta = -0.425642807490658 lketa = 1.62897795656057e-07 wketa = 2.78789813850159e-07 pketa = -1.12422039873405e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.446655722843 lags = 4.24796536201592e-08 wags = -7.35771891609539e-07 pags = -3.081669480013e-14
+ b0 = -1.3225759820552e-07 lb0 = -1.17070457209429e-13 wb0 = 1.29010145139182e-13 pb0 = 1.14195909203109e-19
+ b1 = 5.695485976798e-10 lb1 = -3.24865481301036e-15 wb1 = -5.5556390141237e-16 pb1 = 3.1688873427317e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.139510413282458+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 4.41151957034109e-08 wvoff = 4.62662583074777e-08 pvoff = -3.20031922622566e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '1.57160896883246+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -4.62338504638453e-07 wnfactor = 1.67483167491185e-06 pnfactor = -2.22446162204163e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.98761825507752e-06 lcit = -1.31809774084292e-11 wcit = 3.63621228732703e-12 pcit = 9.56208733703535e-18
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.377419941626962 leta0 = 3.88175157431277e-07 weta0 = 3.33082012678432e-07 peta0 = -3.11685056655008e-13
+ etab = -0.0134909135360391 letab = 2.09302629145866e-08 wetab = 1.26501060949782e-08 petab = -2.06502958804833e-14
+ dsub = -0.0723542883760557 ldsub = 3.24539860205493e-07 wdsub = 2.81697935081916e-07 pdsub = -2.35436143426634e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.28477320981786 lpclm = -4.3051365881767e-06 wpclm = -3.70994057209873e-06 ppclm = 3.12314411734643e-12
+ pdiblc1 = 0.172006588362524 lpdiblc1 = -4.44739713099843e-07 wpdiblc1 = 2.7176167043848e-07 ppdiblc1 = 3.22634645909429e-13
+ pdiblc2 = -0.00342314533019774 lpdiblc2 = 4.89517507092067e-09 wpdiblc2 = 3.95643734416223e-09 ppdiblc2 = -3.55118517449912e-15
+ pdiblcb = -0.025
+ drout = -0.0306258600616882 ldrout = 2.4519821437813e-06 wdrout = 3.31142442250692e-07 pdrout = -1.77878063827757e-12
+ pscbe1 = 398055733.395698 lpscbe1 = 7.68399432421802 wpscbe1 = -86.9948919176757 ppscbe1 = -5.57432294652667e-6
+ pscbe2 = 1.67447714410044e-08 lpscbe2 = -2.36741235002141e-15 wpscbe2 = -1.6183281585089e-15 ppscbe2 = 1.71742981967363e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00211874516120117 lalpha0 = -1.66311362420558e-09 walpha0 = -1.53703512966814e-09 palpha0 = 1.20649912622544e-15
+ alpha1 = -2.901784e-10 walpha1 = 2.830533595664e-16
+ beta0 = 226.361681396106 lbeta0 = -3.65210781637347e-05 wbeta0 = -0.00016203683832208 pbeta0 = 2.64940700695686e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.49173093916349e-07 lagidl = -1.35247964473053e-13 wagidl = -1.08102033897081e-13 pagidl = 9.80768160951437e-20
+ bgidl = 3502305384.9852 lbgidl = -424.017387318792 wbgidl = -1794.61222131597 pbgidl = 0.000307601717560869
+ cgidl = -1649.65663064424 lcgidl = 0.000154985107397515 wcgidl = 0.00285408960760581 pcgidl = -9.63687681278556e-10
+ egidl = 7.85997106636054 legidl = -9.1920358692599e-06 wegidl = -5.04206516207623e-06 pegidl = 6.66832565321111e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.46583137990777 lkt1 = 3.3178676025674e-07 wkt1 = 6.1927400531811e-07 pkt1 = -1.4695893175916e-13
+ kt2 = -0.019032
+ at = -94658.0785163279 lat = 0.113345357890971 wat = 0.097080981749756 pat = -8.82708826559657e-8
+ ute = -1.107123869308 lute = -3.11578271831701e-07 wute = -2.48593028305989e-07 pute = 2.2603321098722e-13
+ ua1 = 2.19843734429792e-09 lua1 = -1.49665945530288e-15 wua1 = -1.19411120727155e-15 pua1 = 1.08574561521166e-21
+ ub1 = 2.29419007058e-18 lub1 = -5.35101814667486e-24 wub1 = -4.26931505134197e-24 pub1 = 3.88187471043269e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.69 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.68355458358111+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.58764448825169e-07 wvth0 = -1.27666416539811e-07 pvth0 = 1.90194453200304e-13
+ k1 = 0.969168697278098 lk1 = -2.42939512574251e-07 wk1 = -2.96945866125607e-07 pk1 = 1.76239497638941e-13
+ k2 = -0.0862168837171923 lk2 = 7.37892120668583e-08 wk2 = 8.09977746140178e-08 pk2 = -4.708947792109e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -143687.962826487 lvsat = 0.110055817862335 wvsat = 0.147107525760443 pvsat = -7.29573108377215e-8
+ ua = -8.40116727511754e-09 lua = 5.59822500444561e-15 wua = 7.56327215925e-15 pua = -4.0568432146054e-21
+ ub = 1.08019103888018e-17 lub = -4.86724806854387e-24 wub = -7.93919264748543e-24 pub = 3.47897315950345e-30
+ uc = -5.14707066768781e-12 luc = 4.17703731275453e-18 wuc = 1.70484682653045e-18 puc = -3.03021501038853e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = -0.00430654062596375 lu0 = 1.28516149780582e-08 wu0 = 1.58689303928379e-08 pu0 = -9.83308699980535e-15
+ a0 = 2.33424232933645 la0 = -9.74359302167535e-07 wa0 = -1.15701551520781e-06 pa0 = 7.0684505832023e-13
+ keta = -0.56219860296167 lketa = 2.87061152688074e-07 wketa = 3.84179228312131e-07 pketa = -2.08247364972953e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 1.05891232734278 lags = 3.95035335978732e-07 wags = -4.54484996317488e-07 pags = -2.86576804344426e-13
+ b0 = -1.18662839188899e-06 lb0 = 8.41616186947265e-13 wb0 = 1.15749191835455e-12 pb0 = -8.20951143092962e-19
+ b1 = -1.365396375285e-08 lb1 = 9.68407379170885e-15 wb1 = 1.33187043268625e-14 pb1 = -9.44629104382723e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0360545754317634+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -4.99520248623329e-08 wvoff = -2.87853654379571e-08 pvoff = 3.623749662828e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '7.27627107179478+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -5.64930252175695e-06 wnfactor = -3.06803649781166e-06 pnfactor = 4.0900067238447e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -7.86924275499999e-05 lcit = 6.29051042398374e-11 wcit = 6.43415667964372e-11 pcit = -4.56342562503731e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.502204453567877 leta0 = -4.11623323899631e-07 weta0 = -3.38125631517002e-07 peta0 = 2.98610493829691e-13
+ etab = 0.0553048603729534 letab = -4.16222945121648e-08 wetab = -4.32696331903175e-08 petab = 3.01947270646719e-14
+ dsub = 0.875511760505652 ldsub = -5.37307344740201e-07 wdsub = -4.05927698615124e-07 pdsub = 3.897874640124e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.14481128275993 lpclm = -1.45012620599927e-06 wpclm = -1.43206775196226e-06 ppclm = 1.05198825563735e-12
+ pdiblc1 = -2.10046491111544 lpdiblc1 = 1.6215049978005e-06 wpdiblc1 = 1.92031702984877e-06 ppdiblc1 = -1.17631431463438e-12
+ pdiblc2 = -0.0615620131490256 lpdiblc2 = 5.77579406351899e-08 wpdiblc2 = 4.61330464478596e-08 ppdiblc2 = -4.1900267002036e-14
+ pdiblcb = -0.025
+ drout = 8.9465792388557 ldrout = -5.71054159240934e-06 wdrout = -6.18133508793853e-06 pdrout = 4.14268955604698e-12
+ pscbe1 = -394403560.362135 lpscbe1 = 728.227607173528 wpscbe1 = 487.891532901768 ppscbe1 = -0.000528289804713607
+ pscbe2 = 2.70650785081174e-08 lpscbe2 = -1.17511515507938e-14 wpscbe2 = -9.10515363911769e-15 ppscbe2 = 8.52482588791718e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000867698582174087 lalpha0 = -5.25599522225207e-10 walpha0 = -6.29468393099262e-10 palpha0 = 3.81294071000188e-16
+ alpha1 = -2.901784e-10 walpha1 = 2.830533595664e-16
+ beta0 = 220.844423845692 lbeta0 = -3.15045117360209e-05 wbeta0 = -0.000158034365901162 pbeta0 = 2.28548220208494e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -5.50465844024042e-08 lagidl = 5.04387780382734e-14 wagidl = 4.00059267095145e-14 pagidl = -3.65903470864038e-20
+ bgidl = -362326022.855995 lbgidl = 3089.89872026082 wbgidl = 1008.96917497679 pbgidl = -0.00224155466701833
+ cgidl = -3552.2174621482 lcgidl = 0.00188488854344249 wcgidl = 0.00329807879980556 pcgidl = -1.36738485428618e-9
+ egidl = -3.10898960757627 legidl = 7.81491623517151e-07 wegidl = 2.91532348298853e-06 pegidl = -5.66929972314023e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.192311711929024 lkt1 = -1.17587984599587e-06 wkt1 = -6.98429728576316e-07 pkt1 = 1.05116318828435e-12
+ kt2 = -0.019032
+ at = -37442.0151 lat = 0.0613216522296749 wat = 0.100377797636235 pat = -9.12685125007462e-8
+ ute = -1.3434125 lute = -9.67328343749982e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.70 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-1.61231625663336+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 3.99959767787138e-07 wvth0 = 6.66164072060669e-07 pvth0 = -3.72829820839586e-13
+ k1 = 0.2061850912346 lk1 = 2.98206610012101e-07 wk1 = 2.36515778323349e-07 pk1 = -2.02118173686482e-13
+ k2 = 0.101930159822552 lk2 = -5.96540785637051e-08 wk2 = -4.61743393372954e-08 pk2 = 4.31073438988788e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -190179.209856701 lvsat = 0.143029734818515 wvsat = 0.204423856067823 pvsat = -1.13608918108231e-7
+ ua = -6.69346222854139e-09 lua = 4.38703520016147e-15 wua = 8.32600612310437e-15 pua = -4.5978122784691e-21
+ ub = 1.74328677397342e-17 lub = -9.57025456969272e-24 wub = -1.62389852089734e-23 pub = 9.36560103373877e-30
+ uc = 8.97113270220401e-12 luc = -5.83629842734124e-18 wuc = -8.44829916268641e-18 puc = 4.17090378246353e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0184673111754759 lu0 = -3.30073941211287e-09 wu0 = 1.30334289984253e-10 pu0 = 1.32951228614358e-15
+ a0 = 1.0278216270047 la0 = -4.77804190387424e-08 wa0 = -3.40371275680225e-07 pa0 = 1.27640131435292e-13
+ keta = -0.58747143159423 lketa = 3.04985906395718e-07 wketa = 4.77397445966158e-07 pketa = -2.74362385844071e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 5.60276787161849 lags = -2.82769420879882e-06 wags = -4.71390934669912e-06 pags = 2.73441991616374e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.375932389042172+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.91106314440849e-07 wvoff = 2.76080561065083e-07 pvoff = -1.79988661744001e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '-10.0362005805755+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 6.62956799768667e-06 wnfactor = 1.12947031968515e-05 pnfactor = -6.09676640459519e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.694333755e-05 lcit = 2.62020621573375e-11 wcit = 3.60362308397973e-11 pcit = -2.55586967231262e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.300492987665518 leta0 = 1.57689836295155e-07 weta0 = 2.72316673646569e-07 peta0 = -1.34345711107572e-13
+ etab = -0.011986611463238 letab = 6.10418188765395e-09 wetab = -2.47130137780409e-09 petab = 1.25851022664674e-15
+ dsub = -0.135768977023096 ldsub = 1.79943518352064e-07 wdsub = 3.74702769896781e-07 pdsub = -1.63874695779669e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.98380930214169 lpclm = -6.2668555124579e-07 wpclm = -6.79558506606253e-07 ppclm = 5.18271073368604e-13
+ pdiblc1 = 1.12885723160216 lpdiblc1 = -6.68891731921964e-07 wpdiblc1 = -5.2011416318386e-07 ppdiblc1 = 5.54561509024015e-13
+ pdiblc2 = 0.0260909508661457 lpdiblc2 = -4.40992409257034e-09 wpdiblc2 = -2.20996885726093e-08 ppdiblc2 = 6.49380031123158e-15
+ pdiblcb = -0.025
+ drout = 4.17525267587675 ldrout = -2.32647822761652e-06 wdrout = -3.77894982228946e-06 pdrout = 2.43879780638538e-12
+ pscbe1 = 1834778071.64029 lpscbe1 = -852.819465324191 wpscbe1 = -1354.36149372574 ppscbe1 = 0.000778328154421953
+ pscbe2 = -9.9097965701732e-10 lpscbe2 = 8.14760770282793e-15 wpscbe2 = 1.13110268664069e-14 ppscbe2 = -5.95535013562613e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000407647910317554 lalpha0 = -1.99308583210961e-10 walpha0 = -3.5902414615968e-10 palpha0 = 1.89481488858288e-16
+ alpha1 = -1.029045151e-09 lalpha1 = 5.2404124314675e-16 walpha1 = 1.00377797636235e-15 palpha1 = -5.11173934462525e-22
+ beta0 = 512.767903388725 lbeta0 = -0.000238551239601917 wbeta0 = -0.000455701668335243 pbeta0 = 2.33975356272221e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.63477859752861e-08 lagidl = -2.85676791521035e-14 wagidl = -9.8518866173956e-14 pagidl = 6.16583622661977e-20
+ bgidl = 11638848237.92 lbgidl = -5421.93412419456 wbgidl = -9012.78693796161 pbgidl = 0.00486637585608324
+ cgidl = -6858.8047645906 lcgidl = 0.00423008558769976 wcgidl = 0.00605529053626084 pcgidl = -3.32293727836709e-9
+ egidl = -12.127467111179 legidl = 7.17784679294738e-06 wegidl = 9.37722191493666e-06 pegidl = -5.15003143517323e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -3.7529476915393 lkt1 = 1.62229538591404e-06 wkt1 = 2.85468488049693e-06 pkt1 = -1.46888334820085e-12
+ kt2 = -0.019032
+ at = 148367.0151 lat = -0.070463402439675 wat = -0.100377797636235 pat = 5.11173934462525e-8
+ ute = -1.83271025 lute = 2.503015948125e-7
+ ua1 = 5.53418499999999e-10 lua1 = -7.22371124999376e-19
+ ub1 = -7.973760125e-18 lub1 = 3.10854354365625e-24
+ uc1 = 4.2331604478072e-10 luc1 = -3.77687004760726e-16 wuc1 = -5.19440645817174e-16 puc1 = 3.68413278045831e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.71 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.096519898550234+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -3.71959527566692e-07 wvth0 = -5.64910762785593e-07 pvth0 = 2.54095038805873e-13
+ k1 = 1.4190614479586 lk1 = -3.19450674649597e-07 wk1 = -5.01293939256023e-07 pk1 = 1.73611424990814e-13
+ k2 = -0.140340584851328 lk2 = 6.3722298161468e-08 wk2 = 7.05856026554891e-08 pk2 = -1.63526565609466e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -456589.290233476 lvsat = 0.278699068250387 wvsat = 0.342101691258066 pvsat = -1.83721355678862e-7
+ ua = 1.15293975258833e-08 lua = -4.89295612977933e-15 wua = -1.04029398198851e-14 pua = 4.93990344299828e-21
+ ub = -2.38981375541509e-17 lub = 1.14775598762183e-23 wub = 2.30065269297307e-23 pub = -1.06201760228963e-29
+ uc = 2.18911233286766e-11 luc = -1.24158036538724e-17 wuc = -1.12835126348696e-17 puc = 5.61473624317284e-24
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.00230154973459434 lu0 = 4.93167460165604e-09 wu0 = 8.74479456460438e-09 pu0 = -3.05740160870673e-15
+ a0 = 1.3516778800476 la0 = -2.12704215900841e-07 wa0 = -1.30421081220629e-08 pa0 = -3.90522471437029e-14
+ keta = -0.37406449461937 lketa = 1.9630842374127e-07 wketa = 1.43021268746883e-07 pketa = -1.04081317595155e-13
+ a1 = 0.0
+ a2 = 0.5
+ ags = 10.1494526938742 lags = -5.14309345453253e-06 wags = -6.77494876233279e-06 pags = 3.78400423857519e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '0.625050838662064+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -3.18644394267533e-07 wvoff = -5.55113653818398e-07 pvoff = 2.43296992185412e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '11.2433570337456+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -4.20704671740637e-06 wnfactor = -6.04282786667115e-06 pnfactor = 2.73237128950374e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 0.0001637269302 lcit = -7.089677169435e-11 wcit = -1.29992255380869e-10 pcit = 5.89913098847482e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.64136744488276 leta0 = 8.40530153633036e-07 weta0 = 1.06540298099835e-06 peta0 = -5.38224913126465e-13
+ etab = 0.122862814740174 letab = -6.25678884064336e-08 wetab = -7.61494695708137e-08 petab = 3.87791173789369e-14
+ dsub = -0.131795651435281 ldsub = 1.77920102296469e-07 wdsub = 3.6823470660901e-07 pdsub = -1.60580834550372e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.94487145956879 lpclm = -2.64385645491554e-06 wpclm = -2.89330393276614e-06 ppclm = 1.64562093164052e-12
+ pdiblc1 = -0.918119203041084 lpdiblc1 = 3.73531017420109e-07 wpdiblc1 = 2.34518477832574e-06 ppdiblc1 = -9.04591976939751e-13
+ pdiblc2 = 0.0995883021168162 lpdiblc2 = -4.18384502169743e-08 wpdiblc2 = -6.64538353427061e-08 ppdiblc2 = 2.90811495539034e-14
+ pdiblcb = 3.168610204 lpdiblcb = -1.626345996387e-06 wpdiblcb = -2.31679174805098e-06 ppdiblcb = 1.17982619769496e-12
+ drout = -6.09480802426281 ldrout = 2.90355018392956e-06 wdrout = 5.14367609384471e-06 pdrout = -2.10504944140595e-12
+ pscbe1 = -7208807731.41374 lpscbe1 = 3752.62660488107 wpscbe1 = 5519.77913352317 ppscbe1 = -0.00272232796000456
+ pscbe2 = 1.60686657065446e-07 lpscbe2 = -7.41867287980867e-14 wpscbe2 = -1.06841693753711e-13 ppscbe2 = 5.42139228401689e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00024980347787622 lalpha0 = -1.18926305990212e-10 walpha0 = -1.12327848364921e-10 palpha0 = 6.38513992063073e-17
+ alpha1 = 0.0
+ beta0 = 171.205652427656 lbeta0 = -6.46106632999923e-05 wbeta0 = -7.97460833266107e-05 pbeta0 = 4.25199746065753e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.12532599970616e-07 lagidl = -3.11804795679225e-13 wagidl = -5.43791072487411e-13 pagidl = 2.88413233331325e-19
+ bgidl = -6435571262.68 lbgidl = 3782.46400648599 wbgidl = 5802.29666508366 pbgidl = -0.00267820546876757
+ cgidl = 12557.44016412 lcgidl = -0.00565763714224611 wcgidl = -0.00864814344750019 pcgidl = 4.16478647786322e-9
+ egidl = 18.8958450671856 legidl = -8.62077493388478e-06 wegidl = -1.29451426890615e-05 pegidl = 6.21763273941286e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.30219587975536 lkt1 = 3.74250025763068e-07 wkt1 = 7.97873602974794e-07 pkt1 = -4.21452205122705e-13
+ kt2 = -0.019032
+ at = 94334.70408 lat = -0.04294744805274 wat = -0.0463358349610197 pat = 2.35965239538993e-8
+ ute = -3.601018991776 lute = 1.15081282156193e-06 wute = 1.72369306054993e-06 pute = -8.77790691085053e-13
+ ua1 = 5.52e-10
+ ub1 = -6.837423648768e-18 lub1 = 2.5298641931351e-24 wub1 = 6.00512421094815e-24 pub1 = -3.05810950442534e-30
+ uc1 = -1.17423208956144e-09 luc1 = 4.35864382653019e-16 wuc1 = 1.03888129163435e-15 puc1 = -4.25162168601357e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.72 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.884106+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.57102
+ k2 = 0.0283423
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 180350.0
+ ua = 2.33445218e-9
+ ub = 9.509e-20
+ uc = -3.2639e-11
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.01916912
+ a0 = 0.87668
+ keta = -0.0076977
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1244
+ b0 = 2.8576e-9
+ b1 = 3.2982e-11
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.10903374+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.5986+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))'
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.99495
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225600350.0
+ pscbe2 = 1.4994384e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.8978653e-5
+ alpha1 = 0.0
+ beta0 = 37.686511
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.74941e-8
+ bgidl = 1701900000.0
+ cgidl = 1200.0
+ egidl = 1.0890786
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.644265
+ kt2 = -0.019032
+ at = 351440.0
+ ute = -1.4104
+ ua1 = 2.2096e-11
+ ub1 = -2.3998e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.73 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.871312129020833+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.54716375791981e-7
+ k1 = 0.561904589374999 lk1 = 1.81480988985786e-7
+ k2 = 0.0303940576565207 lk2 = -4.08489561230881e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 246388.282875 lvsat = -1.3147726833291 wvsat = 4.44089209850063e-16
+ ua = 2.38979930555458e-09 lua = -1.10191975944758e-15
+ ub = -5.45172689583348e-21 lub = 2.00171037620087e-24
+ uc = -2.44202465472083e-11 luc = -1.63629217179993e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0195425091014583 lu0 = -7.43389696820933e-9
+ a0 = 0.857074715876042 la0 = 3.90326502944948e-7
+ keta = -0.00737856176249996 lketa = -6.35380295494683e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.115702210957083 lags = 1.73166456502688e-7
+ b0 = 4.74105606666666e-09 lb0 = -3.74981976952833e-14
+ b1 = 5.4720573625e-11 lb1 = -4.32798696943532e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.109925909991041+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.77624353941467e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.76006074770832+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -3.2145623913121e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.32955208333333e-05 lcit = -6.56113481510418e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.59566989570313 lpclm = -1.19598825835274e-5
+ pdiblc1 = 0.39
+ pdiblc2 = -0.0001257996463375 lpdiblc2 = 2.81875091088449e-08 ppdiblc2 = -2.52435489670724e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 226182167.612082 lpscbe1 = -11.5835522933703
+ pscbe2 = 1.49915241470208e-08 lpscbe2 = 5.6937527925576e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.085503009075e-05 lalpha0 = 5.93966255074515e-10
+ alpha1 = 0.0
+ beta0 = 36.7947648129375 lbeta0 = 1.77539977747748e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.79836769020832e-08 lagidl = -2.08839608937804e-13
+ bgidl = 1821527406.25 lbgidl = -2381.69193788286
+ cgidl = 1068.17916666666 lcgidl = 0.00262445392604166
+ egidl = 0.805099219704164 legidl = 5.65381647715484e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.443169023229165 lkt1 = -4.00367007552473e-6
+ kt2 = -0.019032
+ at = 483491.519791665 lat = -2.62904672041225
+ ute = -1.31436852291666 lute = -1.91191468512132e-6
+ ua1 = 2.2096e-11
+ ub1 = -1.95365238958332e-18 lub1 = -8.88246431268805e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.74 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.922487612937498+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.50043320375922e-7
+ k1 = 0.598366231875001 lk1 = -1.0690325695735e-7
+ k2 = 0.0221870270304375 lk2 = 2.4062500856262e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -17764.8486249996 lvsat = 0.774480471987284
+ ua = 2.16841080333624e-09 lua = 6.49097251722745e-16
+ ub = 3.967151806875e-19 lub = -1.17912823760261e-24
+ uc = -5.72952603583749e-11 luc = 9.63874858059772e-17
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.018048952695625 lu0 = 4.3790140346282e-9
+ a0 = 0.935495852371872 la0 = -2.29925870884749e-7
+ keta = -0.00865511471249999 lketa = 3.74277346484057e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.15049336712875 lags = -1.0200549544807e-7
+ b0 = -2.7927682e-09 lb0 = 2.208870188585e-14
+ b1 = -3.2233720875e-11 lb1 = 2.54944556830594e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.106357230026875+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.04631466124396e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.11421775687501+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 1.89357128393643e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.13437499999977e-07 lcit = 3.8649044453125e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.807209687109375 lpclm = 7.04509275683232e-06 wpclm = 6.35274710440725e-22 ppclm = 1.61558713389263e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00553739893901251 lpdiblc2 = -1.66041443023347e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 223854897.16375 lpscbe1 = 6.82341150011052
+ pscbe2 = 1.50029635589375e-08 lpscbe2 = -3.35396407763159e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00010847970227225 lalpha0 = -3.49881976867543e-10
+ alpha1 = 0.0
+ beta0 = 40.3617495611877 lbeta0 = -1.04581763453225e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.97463070625e-09 lagidl = 1.23019135513408e-13
+ bgidl = 1343017781.25 lbgidl = 1402.96031364845
+ cgidl = 1595.4625 lcgidl = -0.00154596177812499
+ egidl = 1.9410167408875 legidl = -3.33043917726444e-6
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.2475529303125 lkt1 = 2.35840334157415e-6
+ kt2 = -0.019032
+ at = -44714.5593750002 lat = 1.54866721123672
+ ute = -1.69849443125 lute = 1.12623315536405e-6
+ ua1 = 2.2096e-11
+ ub1 = -3.73824283125e-18 lub1 = 5.23230763806401e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.75 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.915353740124999+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 1.22155228083666e-7
+ k1 = 0.5816927075 lk1 = -4.17222817943735e-8
+ k2 = 0.0222051647965 lk2 = 2.39915957942823e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 316049.94375 lvsat = -0.530485005104689
+ ua = 2.6238696406575e-09 lua = -1.13140520807534e-15
+ ub = 4.2981016375e-19 lub = -1.30850480013969e-24 pub = -1.40129846432482e-45
+ uc = -6.11269159088126e-11 luc = 1.11366385266525e-16
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0212460212425001 lu0 = -8.11912618224306e-9
+ a0 = 1.0077881975 la0 = -5.12534721076883e-7
+ keta = 0.0204554322625 lketa = -1.10057632297178e-7
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.16964537764875 lags = 1.14949689257338e-6
+ b0 = -5.80965427249999e-08 lb0 = 2.38284982447707e-13
+ b1 = -3.0793177075e-10 lb1 = 1.33271715830444e-15 wb1 = 1.97215226305253e-31 pb1 = -1.88079096131566e-37
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.14082239165175+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.24269786469604e-7
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.71416690250001+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -4.5177991359814e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0990924999999998 leta0 = -7.46373556250004e-8
+ etab = -0.13682375 letab = 2.61230744687501e-7
+ dsub = 0.792970780341248 ldsub = -9.10741023049034e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.827117569675 lpclm = 6.56098928248008e-7
+ pdiblc1 = 0.240486804332502 lpdiblc1 = 5.84484460163175e-7
+ pdiblc2 = 0.000582952602475005 lpdiblc2 = 2.7640250387746e-9
+ pdiblcb = -0.025
+ drout = 0.68807102942375 ldrout = -5.00661671774797e-7
+ pscbe1 = 175447980.075 lpscbe1 = 196.058152129306
+ pscbe2 = 1.5453002078625e-08 lpscbe2 = -1.79285272386483e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.7096054157625e-05 lalpha0 = -7.08254504754455e-11
+ alpha1 = -9.54625e-11 lalpha1 = 3.73186778125001e-16
+ beta0 = 70.7991215633749 lbeta0 = -0.000129445472844874
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.3615720574875e-08 lagidl = -1.0211594523233e-13
+ bgidl = 2344744475.0 lbgidl = -2513.03976389374
+ cgidl = 751.326250000006 lcgidl = 0.00175397785718749
+ egidl = 1.2603426589975 legidl = -6.69514022635976e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.739493616875002 lkt1 = 3.72272470518589e-7
+ kt2 = -0.019032
+ at = 653712.460000001 lat = -1.181658614255
+ ute = -1.372787775 lute = -1.47035590581247e-7
+ ua1 = -4.84145456e-10 lua1 = 1.979024411868e-15 wua1 = -1.97215226305253e-31 pua1 = 1.22251412485518e-36
+ ub1 = -1.2627461625e-18 lub1 = -4.44502771424685e-24
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.76 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.847360479749998+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -7.66090428730976e-9
+ k1 = 0.55984
+ k2 = 0.0343814394499999 lk2 = 7.44043412087399e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9715.01600000006 lvsat = 0.054384955702
+ ua = 2.03140494945e-09 lua = -2.41996387415246e-19
+ ub = -2.87190992499999e-19 lub = 6.04296574306256e-26
+ uc = -2.7970035e-12
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0171738952000001 lu0 = -3.44419535600007e-10
+ a0 = 0.73934
+ keta = -0.0413415447499998 lketa = 7.92824606393747e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.43242187
+ b0 = 4.557803e-08 lb0 = 4.03443044725e-14
+ b1 = -1.96275324999999e-10 lb1 = 1.11953708925626e-15 pb1 = -7.52316384526264e-37
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.075734118+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.88030138000002+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -7.68972164764994e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08172107325 leta0 = -4.14709591025627e-8
+ etab = 0.003946781475 letab = -7.53539253114375e-9
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.1707598
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 278136550.0
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.58509926525e-10 lagidl = -5.27658019678568e-17
+ bgidl = 1028500000.0
+ cgidl = 2284.598445 lcgidl = -0.00117342208111626
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.612185477499999 lkt1 = 1.29209405416875e-7
+ kt2 = -0.019032
+ at = 39164.4 lat = -0.00833273069999996
+ ute = -1.4498
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.77 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.859537932499997+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 3.41144462562981e-9
+ k1 = 0.55984
+ k2 = 0.0254354992500003 lk2 = 8.87813953893724e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 59094.2232499998 lvsat = 0.00948691150993719
+ ua = 2.02451866050001e-09 lua = 6.01936184037006e-18
+ ub = -1.41967787499997e-19 lub = -7.16145417156231e-26
+ uc = -2.7970035e-12
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0175681825 lu0 = -7.02925263125037e-10
+ a0 = 0.73934
+ keta = -0.032622
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.43242187
+ b0 = 4.0893064125e-07 lb0 = -2.90034057306562e-13
+ b1 = 4.70536875e-09 lb1 = -3.3372827859375e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.075734118+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))'
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.04709826249999+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.13822301781019e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.036111
+ etab = -0.0043407
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.1707598
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 278136550.0
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.00079456125001e-10 lagidl = 3.62103243344307e-19
+ bgidl = 1028500000.0
+ cgidl = 994.06
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.770447375000003 lkt1 = 2.7310903571875e-7
+ kt2 = -0.019032
+ at = 100925.0 lat = -0.0644885562499999
+ ute = -1.34341249999999 lute = -9.67328343749914e-8
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.78 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.69403416250001+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.13972104246875e-7
+ k1 = 0.532213187500002 lk1 = 1.95943167656254e-8
+ k2 = 0.0382805713799999 lk2 = -2.32227869265155e-10
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 91611.3797499994 lvsat = -0.0135758817376876
+ ua = 4.78362376146251e-09 lua = -1.95087593101728e-15
+ ub = -4.95196201875e-18 lub = 3.33987386679844e-24 pub = -1.40129846432482e-45
+ uc = -2.67452963887499e-12 luc = -8.68645860029027e-20
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0186469720875 lu0 = -1.46805677805944e-9
+ a0 = 0.558632637499997 la0 = 1.28166696853125e-7
+ keta = 0.0706029749999999 lketa = -7.32123135187498e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.895178697387497 lags = 9.41600702419583e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '0.00463427073+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -5.70012797067521e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.53312256249998+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.77459496495313e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.273125e-05 lcit = -9.02963906250003e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.0748852950000003 leta0 = -2.75006687287499e-8
+ etab = -0.015393207375 letab = 7.83899085571874e-9
+ dsub = 0.380744684775001 ldsub = -4.59515803591676e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.04706348425 lpclm = 8.7731611945689e-8
+ pdiblc1 = 0.411899438487506 lpdiblc1 = 9.5550430587743e-8
+ pdiblc2 = -0.00437263784012498 lpdiblc2 = 4.54153516315867e-9
+ pdiblcb = -0.025
+ drout = -1.03388738732501 ldrout = 1.03531273461276e-6
+ pscbe1 = -32158259.5625 lpscbe1 = 220.076593682203
+ pscbe2 = 1.46008450500001e-08 lpscbe2 = -6.16182569624666e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -8.7253358915e-05 lalpha0 = 6.18845157354639e-11 walpha0 = -2.90265314380597e-26 palpha0 = -3.29574761733266e-32
+ alpha1 = 3.54625e-10 lalpha1 = -1.8059278125e-16
+ beta0 = -115.39969052625 lbeta0 = 8.39749805057428e-05 wbeta0 = 6.7762635780344e-20 pbeta0 = -2.58493941422821e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.94567620874998e-08 lagidl = 5.64260519680593e-14 wagidl = 7.49417859959961e-30 pagidl = -2.82118644197349e-35
+ bgidl = -784939250.0 lbgidl = 1286.1817880625
+ cgidl = 1488.185275 lcgidl = -0.000350458351293749
+ egidl = 0.798680272550001 legidl = 7.8722343748911e-8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.182127945375001 lkt1 = -4.0250501025722e-7
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.83271025000001 lute = 2.50301594812498e-7
+ ua1 = 5.53418500000001e-10 lua1 = -7.22371125001742e-19
+ ub1 = -7.97376012499999e-18 lub1 = 3.10854354365625e-24
+ uc1 = -2.9271333e-10 luc1 = 1.301568293025e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.79 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 7e-07 wmax = 7.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.875228117749984+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.16990825358093e-8
+ k1 = 0.728046624999998 lk1 = -8.01338612812541e-8
+ k2 = -0.0430409889400005 lk2 = 4.11807767236951e-8
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 14985.0120000001 lvsat = 0.0254460960389999
+ ua = -2.81066337442502e-09 lua = 1.91651479293344e-15
+ ub = 7.8154936875e-18 lub = -3.16195295160938e-24 pub = -5.60519385729927e-45
+ uc = 6.33722595400001e-12 luc = -4.67610112167453e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0143559198249998 lu0 = 7.1716158661875e-10
+ a0 = 1.333699825 la0 = -2.66536268381248e-7
+ keta = -0.17691506 lketa = 5.2836245805e-8
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.810440882749987 lags = 7.3013931234561e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.140152434659999+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.67313500131051e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.91354631499999+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -4.40575760913748e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.54625000000001e-05 lcit = 1.0420528125e-11
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.172749545000001 leta0 = 9.86073735412505e-8
+ etab = 0.01789363775 letab = -9.11233502418751e-9
+ dsub = 0.375802028624996 ldsub = -4.34345327147821e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.95656091299999 lpclm = -3.75429953645253e-7
+ pdiblc1 = 2.314629724275 lpdiblc1 = -8.73414967449549e-07 ppdiblc1 = 1.61558713389263e-27
+ pdiblc2 = 0.00798419189674998 lpdiblc2 = -1.75118038034497e-9
+ pdiblcb = -0.025
+ drout = 0.995555826174993 ldrout = 1.81877813788242e-9
+ pscbe1 = 400000000.0
+ pscbe2 = 1.34094045149998e-08 lpscbe2 = 5.45122835486235e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.49637677324995e-05 lalpha0 = -3.09095560097756e-11
+ alpha1 = 0.0
+ beta0 = 61.2786787774994 lbeta0 = -5.99847906219216e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.3706292125e-07 lagidl = 8.57619885215628e-14
+ bgidl = 1562676249.99998 lbgidl = 90.6585946875057
+ cgidl = 636.300000000003 lcgidl = 8.33642250000037e-5
+ egidl = 1.05145321849999 legidl = -5.00022789761254e-8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.202357155749993 lkt1 = -2.06705972509311e-7
+ kt2 = -0.019032
+ at = 30462.5000000001 lat = -0.0104205281250001
+ ute = -1.22497299999999 lute = -5.91885997499944e-8
+ ua1 = 5.52e-10
+ ub1 = 1.44041400000003e-18 lub1 = -1.68562462950001e-24
+ uc1 = 2.57826660000001e-10 luc1 = -1.50205660605e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.80 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.840842795292857+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0 = -2.92219585666209e-8
+ k1 = 0.526122755928571 wk1 = 3.03256639190702e-8
+ k2 = 0.0374742384411143 wk2 = -6.16813129229688e-9
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 397324.158664286 wvsat = -0.146554327573157
+ ua = 3.39404775977e-09 wua = -7.15699595973328e-16
+ ub = -1.00436427687857e-18 wub = 7.42621993500524e-25
+ uc = -1.98255285019357e-11 wuc = -8.65480806948153e-18
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0203424788973571 wu0 = -7.92540573784292e-10
+ a0 = 0.837601461357143 wa0 = 2.63954426121635e-8
+ keta = -0.0126323011571429 wketa = 3.33305661318751e-9
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.1478249358405 wags = -1.58222792137223e-8
+ b0 = 3.13121993914286e-08 wb0 = -1.92195453405429e-14
+ b1 = -1.5890781751e-09 wb1 = 1.09561405703059e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0904679739921428+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' wvoff = -1.25401723869431e-8
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.31416134142857+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor = 1.92122954177438e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.39933134797885e-05 wcit = -9.45172761666919e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.28215321075893 wpclm = -8.69436259894275e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 226448228.593214 wpscbe1 = -0.572696204272233
+ pscbe2 = 1.49864524830857e-08 wpscbe2 = 5.35731137369028e-18
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.57821989629929e-05 walpha0 = -1.81043479065197e-11
+ alpha1 = -1.41230714285714e-10 walpha1 = 9.53937210414286e-17
+ beta0 = 86.6745182460929 wbeta0 = -3.30887535423444e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.12219718014286e-08 wagidl = -2.27813560967877e-14
+ bgidl = 2345347134.28571 wbgidl = -434.613793064749
+ cgidl = 917.538571428571 wcgidl = 0.000190787442082857
+ egidl = -0.197422199801429 wegidl = 8.68961819222676e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.133765398607143 wkt1 = -3.448149137624e-7
+ kt2 = -0.019032
+ at = 781685.248 wat = -0.290607431780608
+ ute = -1.36181663428571 wute = -3.28154400382512e-8
+ ua1 = -9.44577396228572e-10 wua1 = 6.52935678789004e-16
+ ub1 = -1.34734871714286e-18 wub1 = -7.10874009200726e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.81 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.827684028164882+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.61981184442637e-07 wvth0 = -2.94684262107489e-08 pvth0 = 4.90698594385608e-15
+ k1 = 0.459936470600921 lk1 = 1.31771930115953e-06 wk1 = 6.88739579534765e-08 pk1 = -7.67467623004505e-13
+ k2 = 0.0539776717677458 lk2 = -3.28570979958239e-07 wk2 = -1.59294578169705e-08 pk2 = 1.94340690111357e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 606371.013573911 lvsat = -4.16196609610946 wvsat = -0.243148895519657 pvsat = 1.92312540188885e-6
+ ua = 4.11353301065253e-09 lua = -1.43244117311331e-14 wua = -1.16428903617359e-15 pua = 8.93107931230704e-21
+ ub = -1.79193843023888e-18 lub = 1.56800107127887e-23 wub = 1.20667529782625e-24 pub = -9.23895324914691e-30
+ uc = 9.46346888351422e-12 luc = -5.83121971196268e-16 wuc = -2.28866200528198e-17 puc = 2.83344702729277e-22
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0230700625245941 lu0 = -5.43041443305667e-08 wu0 = -2.38267184944333e-09 pu0 = 3.16583210999148e-14
+ a0 = 0.767641113755024 la0 = 1.39285805049748e-06 wa0 = 6.04075688182328e-08 pa0 = -6.77155923668189e-13
+ keta = -0.0127459185818393 lketa = 2.26203771263703e-09 wketa = 3.62535969419543e-09 pketa = -5.81953511555689e-15
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.137358433727713 lags = 2.08380207189007e-07 wags = -1.46276090455306e-08 pags = -2.37849870460713e-14
+ b0 = 5.7556755335655e-08 lb0 = -5.22509425432588e-13 wb0 = -3.5674152808441e-14 pb0 = 3.27598893730251e-19
+ b1 = -2.21717868477166e-09 lb1 = 1.25050100721804e-14 wb1 = 1.53454526648699e-15 pb1 = -8.73879118186966e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.0972535891294481+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.35096508172395e-07 wvoff = -8.55946843667992e-09 pvoff = -7.92528301217766e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.29780037661942+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 3.25734538626708e-07 wnfactor = 3.12231918610526e-07 pnfactor = -2.39127940013946e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.41847417269476e-05 lcit = -2.02903692829753e-10 wcit = -1.41095406957082e-11 pcit = 9.2733565043857e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.7312738733056 lpclm = -2.88509055508072e-05 wpclm = -1.44248516425568e-06 ppclm = 1.14089738991573e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00192601428407009 lpdiblc2 = -1.26625673851222e-08 wpdiblc2 = -1.38588951203808e-09 ppdiblc2 = 2.75920207675441e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 227851751.374683 lpscbe1 = -27.9430859369559 wpscbe1 = -1.1277136741129 ppscbe1 = 1.10499815614254e-5
+ pscbe2 = 1.49795536393166e-08 lpscbe2 = 1.3735080531124e-16 wpscbe2 = 8.08543154682739e-18 ppscbe2 = -5.43148265571155e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.61858078545599e-05 lalpha0 = 1.43282903973236e-09 walpha0 = 1.03551125174543e-11 palpha0 = -5.66606512446003e-16
+ alpha1 = -1.41230714285714e-10 walpha1 = 9.53937210414286e-17
+ beta0 = 84.5233525494264 lbeta0 = 4.28280956463573e-05 wbeta0 = -3.22380836722605e-05 pbeta0 = -1.69361991109694e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.37935370230555e-08 lagidl = -6.48475434888674e-13 wagidl = -3.76965467792701e-14 pagidl = 2.96950260095212e-19
+ bgidl = 2683912229.82072 lbgidl = -6740.5771282802 wbgidl = -582.494379541545 pbgidl = 0.00294419156631316
+ cgidl = 678.669123011161 lcgidl = 0.00475571156590434 wcgidl = 0.000263093000946937 pcgidl = -1.43954944781468e-9
+ egidl = -0.882467687313214 legidl = 1.3638741872244e-05 wegidl = 1.13986031707726e-06 pegidl = -5.3933859184114e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.401485157292445 lkt1 = -1.06564371300439e-05 wkt1 = -5.705182876166e-07 pkt1 = 4.49358489590674e-12
+ kt2 = -0.019032
+ at = 1197313.203437 lat = -8.2748408717841 wat = -0.482148000931506 pat = 3.81342907636752e-6
+ ute = -1.2337636584294 lute = -2.54943870956723e-06 wute = -5.44442332984628e-08 pute = 4.3061305221587e-13
+ ua1 = -1.58171585948864e-09 lua1 = 1.26849489496605e-14 wua1 = 1.08328830524417e-15 pua1 = -8.56799802825242e-21
+ ub1 = -2.07526080981368e-19 lub1 = -2.26930138189981e-23 wub1 = -1.17941403063996e-24 pub1 = 9.32828042183913e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.82 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.93968596890534+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 6.2387016535884e-07 wvth0 = 1.16165607450544e-08 pvth0 = -3.2004444713633e-13
+ k1 = 0.707649136572531 lk1 = -6.41502102176437e-07 wk1 = -7.38147008463289e-08 pk1 = 3.61092651607855e-13
+ k2 = -0.0132742576234499 lk2 = 2.03341342579076e-07 wk2 = 2.39521828743296e-08 pk2 = -1.21093176526308e-13
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -100746.405949161 lvsat = 1.4308023542534 wvsat = 0.0560495609683751 pvsat = -4.43309990089121e-7
+ ua = 1.96898556424438e-09 lua = 2.63735015937067e-15 wua = 1.34700980043648e-16 pua = -1.34295747345914e-21
+ ub = 9.07325468770689e-19 lub = -5.66914228045273e-24 wub = -3.44889676644638e-25 pub = 3.03276202518694e-30
+ uc = -8.8016583062436e-11 luc = 1.87872129657239e-16 wuc = 2.07505945351672e-17 puc = -6.1792936750759e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.015611385368136 lu0 = 4.68839796914935e-09 wu0 = 1.64644510108313e-09 pu0 = -2.08972141036682e-16
+ a0 = 0.91725446135687 la0 = 2.09528680977588e-07 wa0 = 1.23210745955212e-08 pa0 = -2.96827819237209e-13
+ keta = -0.0134730941130139 lketa = 8.01345078258025e-09 wketa = 3.25428491415953e-09 pketa = -2.88461191155795e-15
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.188921082839435 lags = -1.99441675297882e-07 wags = -2.59558468659194e-08 pags = 6.58128779348392e-14
+ b0 = -5.59252475015429e-09 lb0 = -2.30459819139011e-14 wb0 = 1.89108436277551e-15 pb0 = 3.04860416338067e-20
+ b1 = 7.87936778220946e-09 lb1 = -6.73511000717901e-14 wb1 = -5.34385958885239e-15 pb1 = 4.56642324202233e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.103294200073153+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 1.82873210278897e-07 wvoff = -2.06891133012141e-09 pvoff = -1.30588268916825e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.15937673256042+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 9.32981174540034e-06 wnfactor = 6.44943550509189e-07 pnfactor = -5.02277887473398e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.93541795758929e-07 lcit = 6.59412052260009e-11 wcit = -5.41061261531853e-14 pcit = -1.84343808253959e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.391512794734925 lpclm = 3.75724490339227e-06 wpclm = -2.80780803166753e-07 ppclm = 2.22076368121467e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -0.000618042852210232 lpdiblc2 = 7.45901652000288e-09 wpdiblc2 = 4.15766853611423e-09 ppdiblc2 = -1.62533657248046e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 222239647.83102 lpscbe1 = 16.4444440157649 wpscbe1 = 1.09101370079549 ppscbe1 = -6.49848792856839e-6
+ pscbe2 = 1.50071641973129e-08 lpscbe2 = -8.10280005212059e-17 wpscbe2 = -2.83730438809909e-18 ppscbe2 = 3.20758226362267e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000292135247352967 lalpha0 = -1.08485176616777e-09 walpha0 = -1.2404940330259e-10 palpha0 = 4.96432404303683e-16
+ alpha1 = -2.79257256741071e-10 lalpha1 = 1.09168643091503e-15 walpha1 = 1.8862319703673e-16 palpha1 = -7.37375233015836e-22
+ beta0 = 140.006817433176 lbeta0 = -0.000396004498985439 wbeta0 = -6.73048625138631e-05 pbeta0 = 2.60415721441977e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.09201552640111e-08 lagidl = 2.58823835832807e-13 wagidl = 1.14457867804415e-14 pagidl = -9.1728741611937e-20
+ bgidl = 1798581290.64695 lbgidl = 261.726602379891 wbgidl = -307.708550168132 pbgidl = 0.000770841745341491
+ cgidl = 1358.09383177009 lcgidl = -0.000618028311847221 wcgidl = 0.00016032971748122 pcgidl = -6.26768948063461e-10
+ egidl = 0.931783768626985 legidl = -7.10626455651027e-07 wegidl = 6.81682374181476e-07 pegidl = -1.76954202356291e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -1.61812272221642 lkt1 = 5.31714649096162e-06 wkt1 = 2.50299883662333e-07 pkt1 = -1.99847122528117e-12
+ kt2 = -0.019032
+ at = -226619.739676915 lat = 2.98740075853964 wat = 0.122867126414207 pat = -9.7178681959157e-7
+ ute = -1.74266292483571 lute = 1.47557281325687e-06 wute = 2.98334323184961e-08 pute = -2.35960074565065e-13
+ ua1 = 2.2096e-11
+ ub1 = -3.73824283125e-18 lub1 = 5.23230763806406e-24 wub1 = 7.3468396926393e-40
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.83 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.866503364593246+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 3.37781069451782e-07 wvth0 = -3.29957907514206e-08 pvth0 = -1.45643612048735e-13
+ k1 = 0.570536840417053 lk1 = -1.05495858430633e-07 wk1 = 7.53518579770808e-09 pk1 = 4.30756072446547e-14
+ k2 = 0.0211236485151043 lk2 = 6.88713280069334e-08 wk2 = 7.30505846203609e-10 pk2 = -3.03138356041063e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 606925.984782384 lvsat = -1.33566593921389 wvsat = -0.19647105841116 pvsat = 5.43856241220326e-7
+ ua = 3.130492997952e-09 lua = -1.90327277585086e-15 wua = -3.42196720191142e-16 pua = 5.21354861183709e-22
+ ub = 4.48162819360829e-19 lub = -3.87416069324723e-24 wub = -1.23962278217115e-26 pub = 1.73296201037592e-30
+ uc = -8.71629883022944e-11 luc = 1.84535214341155e-16 wuc = 1.75859609538878e-17 puc = -4.94215929231423e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0216594220214879 lu0 = -1.89548893179665e-08 wu0 = -2.79229902564238e-10 pu0 = 7.31897286697178e-15
+ a0 = 1.38150154103959 la0 = -1.60532921527209e-06 wa0 = -2.52423183040441e-07 pa0 = 7.38123669926179e-13
+ keta = 0.0511785059911215 lketa = -2.44725816924511e-07 wketa = -2.07517772577025e-08 pketa = 9.09610866337937e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = -0.591430739362616 lags = 2.85114868564549e-06 wags = 2.84893235428184e-07 pags = -1.14937389702339e-12
+ b0 = -1.90440337582046e-07 lb0 = 6.99570330399172e-13 wb0 = 8.93910868610123e-14 pb0 = -3.11573343132425e-19
+ b1 = -9.94368632850886e-09 lb1 = 2.32367421053554e-15 wb1 = 6.50843187301999e-15 pb1 = -6.69337977101286e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.128678481183172+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 2.82106711208236e-07 wvoff = -8.2025557503591e-09 pvoff = -1.0661031946701e-13
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '4.18057720896095+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 1.42843378303157e-06 wnfactor = -3.15034975857821e-07 pnfactor = -1.26998282053374e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.70615357142857e-05 wcit = -4.76968605207143e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.678828693687501 leta0 = -2.34097107079786e-06 weta0 = -3.91580493081447e-07 peta0 = 1.53078604257865e-12
+ etab = -1.56122209565313 letab = 5.82955997743198e-06 wetab = 9.62104164978021e-07 petab = -3.76110570694033e-12
+ dsub = 0.7175299656192 ldsub = -6.15824018096858e-07 wdsub = 5.09561965407498e-08 pdsub = -1.99200511326927e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.942230264434945 lpclm = -1.45669015066754e-06 wpclm = -7.77524092248252e-08 ppclm = 1.42707493219719e-12
+ pdiblc1 = 0.290083303113651 lpdiblc1 = 3.9059934730296e-07 wpdiblc1 = -3.34997567157334e-08 ppdiblc1 = 1.3095892394098e-13
+ pdiblc2 = -0.000415615487388112 lpdiblc2 = 6.66767734407198e-09 wpdiblc2 = 6.7447882202568e-10 ppdiblc2 = -2.63670633500389e-15
+ pdiblcb = -0.025
+ drout = 0.532271120345961 ldrout = 1.08399122787553e-07 wdrout = 1.05234425386957e-07 pdrout = -4.11387677443959e-13
+ pscbe1 = 196925193.479901 lpscbe1 = 115.404974687874 wpscbe1 = -14.5066978854868 ppscbe1 = 5.44768660901051e-5
+ pscbe2 = 1.57444833774769e-08 lpscbe2 = -2.96339300557747e-15 wpscbe2 = -1.96879877384328e-16 ppscbe2 = 7.90636751121704e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.63671642285064e-05 lalpha0 = -8.49903872134746e-11 walpha0 = 4.92325787063427e-13 palpha0 = 9.56764985995477e-18
+ alpha1 = -2.30284870625e-10 lalpha1 = 9.00241130490782e-16 walpha1 = 9.10652309491738e-17 palpha1 = -3.55996754088058e-22
+ beta0 = 116.302829182779 lbeta0 = -0.000303339682917574 wbeta0 = -3.07352972966958e-05 pbeta0 = 1.17456148616765e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.22898488886915e-07 lagidl = -3.03399198814202e-13 wagidl = -4.67967687252944e-14 pagidl = 1.35955968498861e-19
+ bgidl = 3393232968.29911 lbgidl = -5972.16546848183 wbgidl = -708.197358844914 pbgidl = 0.0023364526206612
+ cgidl = 52.9463701624991 lcgidl = 0.00448411940244225 wcgidl = 0.00047171789631672 pcgidl = -1.84406318617614e-9
+ egidl = 1.36123605950939 legidl = -2.38946282378308e-06 wegidl = -6.81480438021556e-08 pegidl = 1.1617325379396e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.445040686447647 lkt1 = 7.31275542632545e-07 wkt1 = -1.98887054045434e-07 pkt1 = -2.4248718904708e-13
+ kt2 = -0.019032
+ at = 1218677.79757633 lat = -2.66262863896761 wat = -0.381603577404582 pat = 1.00031527931203e-6
+ ute = -1.14989806194482 lute = -8.41693226999349e-07 wute = -1.50549965124268e-07 pute = 4.69203721888059e-13
+ ua1 = -4.84145456e-10 lua1 = 1.979024411868e-15 wua1 = 1.23259516440783e-32 pua1 = 1.6456920911512e-37
+ ub1 = -7.40579121069375e-19 lub1 = -6.48630922095955e-24 wub1 = -3.5269563946615e-25 pub1 = 1.37877542858305e-30
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.84 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.624983659588368+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.23340427328783e-07 wvth0 = -1.50203533670894e-07 pvth0 = 7.81352711202689e-14
+ k1 = 0.503704709980127 lk1 = 2.21033866060673e-08 wk1 = 3.79163571027631e-08 pk1 = -1.49296440695218e-14
+ k2 = 0.0642352303839229 lk2 = -1.34394596761085e-08 wk2 = -2.01646236711545e-08 pk2 = 9.58019042690965e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -214379.234045022 lvsat = 0.232411049832332 wvsat = 0.15136356481591 pvsat = -1.20247013175956e-7
+ ua = 1.87853865551165e-09 lua = 4.87021052453392e-16 wua = 1.03252926775485e-16 pua = -3.29119877287325e-22
+ ub = -2.25827341519289e-18 lub = 1.29310268757446e-24 wub = 1.33135973807822e-24 pub = -8.32604067518531e-31
+ uc = 1.87376118191254e-11 luc = -1.76555064406657e-17 wuc = -1.45454697788419e-17 puc = 1.19253412033219e-23
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0090222293922905 lu0 = 5.1726707093286e-09 wu0 = 5.50601006315415e-09 pu0 = -3.72649653757605e-15
+ a0 = 0.223987006477121 la0 = 6.04655409841307e-07 wa0 = 3.48093118063055e-07 pa0 = -4.08412077955671e-13
+ keta = -0.0916345537048743 lketa = 2.79400173000688e-08 wketa = 3.3970211726534e-08 pketa = -1.35168708343599e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 0.938020096526634 lags = -6.89553227760645e-08 wags = -3.41504299714509e-07 pags = 4.65755969478017e-14
+ b0 = 1.13084654792293e-07 lb0 = 1.20065238708465e-13 wb0 = -4.5597079689455e-14 pb0 = -5.38471861459456e-20
+ b1 = 4.90008365631265e-08 lb1 = -1.10216156120319e-13 wb1 = -3.32299924363875e-14 pb1 = 7.52012486356349e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '0.0777396112438548+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.11997031758065e-07 wvoff = -1.03663216522845e-07 pvoff = 7.56479471128578e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '5.8338848178611+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -1.72814376926107e-06 wnfactor = -1.31954011876953e-06 pnfactor = 6.47868623570452e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.70615357142857e-05 wcit = -4.76968605207143e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -0.755009624295931 leta0 = 3.96584737812006e-07 weta0 = 5.65166402734609e-07 peta0 = -2.95882968258157e-13
+ etab = 2.85732551640859 letab = -2.60655205089684e-06 wetab = -1.92730325299595e-06 petab = 1.75549540582648e-12
+ dsub = 0.405659522968226 ldsub = -2.03853754654855e-08 wdsub = -6.05900816541365e-08 pdsub = 1.37692203166602e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.976434170096058 lpclm = 2.20651992096078e-06 wpclm = 1.4503135783255e-06 ppclm = -1.49038505453327e-12
+ pdiblc1 = 0.285578880888783 lpdiblc1 = 3.9919941543579e-07 wpdiblc1 = 1.76319058158915e-07 ppdiblc1 = -2.69637648358442e-13
+ pdiblc2 = 0.00292590661234337 lpdiblc2 = 2.8787627515964e-10 wpdiblc2 = -6.04694390729282e-10 ppdiblc2 = -1.94444878551478e-16
+ pdiblcb = -0.025
+ drout = 1.31540614772142 ldrout = -1.38680142822903e-06 wdrout = -6.00852862781459e-07 pdrout = 9.36709477491588e-13
+ pscbe1 = 278095801.623538 lpscbe1 = -39.5700089103636 wpscbe1 = 0.0275233278881046 ppscbe1 = 2.67274042384695e-5
+ pscbe2 = 1.43747816404678e-08 lpscbe2 = -3.48289964192794e-16 wpscbe2 = 9.40121943545987e-17 ppscbe2 = 2.35251063154164e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.02943896600239e-06 lalpha0 = -1.16816725643586e-11 walpha0 = 1.37084397643045e-12 palpha0 = 7.89033900690577e-18
+ alpha1 = 2.41230714285714e-10 walpha1 = -9.53937210414286e-17
+ beta0 = -36.2326700435501 lbeta0 = -1.21112810197054e-05 wbeta0 = 2.64995500502357e-05 pbeta0 = 8.18051631963596e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -4.91742027584622e-08 lagidl = 2.5130587709735e-14 wagidl = 3.33215834522238e-14 pagidl = -1.70099953960656e-20
+ bgidl = 542491006.726049 lbgidl = -529.386378348453 wbgidl = 328.272830470918 pbgidl = 0.000357571911709949
+ cgidl = 3688.98599787668 lcgidl = -0.00245798925677105 wcgidl = -0.000948587955040342 pcgidl = 8.67655760527332e-10
+ egidl = -0.805065380093374 legidl = 1.74654819977851e-06 wegidl = 1.15821389585331e-06 pegidl = -1.17969899534759e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.0309563063917961 lkt1 = -5.93150599890881e-08 wkt1 = -3.92588918708352e-07 pkt1 = 1.27338096060596e-13
+ kt2 = -0.019032
+ at = -388828.359337858 lat = 0.406502491120804 wat = 0.289085997323718 pat = -2.80198791237975e-7
+ ute = -1.7189054517675 lute = 2.44684132019599e-07 wute = 1.81766200974551e-07 pute = -1.6527091823611e-13
+ ua1 = 5.524e-10
+ ub1 = -3.74275659545947e-18 lub1 = -7.54401877980269e-25 wub1 = 1.02570929976714e-25 pub1 = 5.0955773087426e-31
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.85 pmos
* DC IV MOS Parameters
+ lmin = 8.0e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.811016126094035+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = 4.58095928414947e-08 wvth0 = -3.2773860049684e-08 pvth0 = -2.86376596198161e-14
+ k1 = 0.243980432776477 lk1 = 2.58257685653486e-07 wk1 = 2.13346081242859e-07 pk1 = -1.74439120743904e-13
+ k2 = 0.119077892628627 lk2 = -6.33051503221058e-08 wk2 = -6.32503800380201e-08 pk2 = 4.87559144034822e-14
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -50339.2695440225 lvsat = 0.0832577121097989 wvsat = 0.0739164149737513 pvsat = -4.98281921819741e-8
+ ua = 1.42235618029067e-09 lua = 9.01804968048055e-16 wua = 4.06728238607467e-16 pua = -6.05054804570556e-22
+ ub = 1.32430037293605e-18 lub = -1.96435252928178e-24 wub = -9.90384963893887e-25 pub = 1.27844230274961e-30
+ uc = -9.77788698200028e-13 luc = 2.7072147971244e-19 wuc = -1.22878136101658e-18 puc = -1.82857740585849e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.016015799993073 lu0 = -1.18623335943289e-09 wu0 = 1.0485505547738e-09 pu0 = 3.26448520418783e-16
+ a0 = 1.54962366890774 la0 = -6.0067972547373e-07 wa0 = -5.47302863029054e-07 pa0 = 4.05726717852329e-13
+ keta = -0.146203127647765 lketa = 7.75564931576423e-08 wketa = 7.67179183451723e-08 pketa = -5.23852230773568e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = 2.25366146975215 lags = -1.26520224138137e-06 wags = -1.23014900269419e-06 pags = 8.5457579313208e-13
+ b0 = 1.11443730539179e-06 lb0 = -7.90414658849124e-13 wb0 = -4.76531654267912e-13 pb0 = 3.37980075789517e-19
+ b1 = -3.28310727376482e-07 lb1 = 2.3285438339177e-13 wb1 = 2.24934390064248e-13 pb1 = -1.59534716153068e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.109982260050812+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = 5.86890797166114e-08 wvoff = 2.3132770555653e-08 pvoff = -3.96413041382663e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '2.74294756778051+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = 1.08229092537471e-06 wnfactor = 2.05437370145501e-07 pnfactor = -7.38717158225544e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.70615357142857e-05 wcit = -4.76968605207143e-12
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.695657588329999 leta0 = -9.22434425268122e-07 weta0 = -4.45488104901144e-07 peta0 = 6.23054642809652e-13
+ etab = -0.00554228387326099 letab = -3.4895034905717e-09 wetab = 8.1160502085864e-10 petab = 2.35697117469269e-15
+ dsub = 1.38934213887555 ldsub = -9.14798793979221e-07 wdsub = -7.25014569838275e-07 pdsub = 6.17897186198088e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.56027446049933 lpclm = -9.99824014080783e-08 wpclm = -2.63096119375627e-07 ppclm = 6.75327131014804e-14
+ pdiblc1 = 0.629864740670508 lpdiblc1 = 8.61574974292555e-08 wpdiblc1 = -5.62274486872123e-08 ppdiblc1 = -5.81947370086009e-14
+ pdiblc2 = 0.0298828119730369 lpdiblc2 = -2.4222689924051e-08 wpdiblc2 = -1.88126282889883e-08 ppdiblc2 = 1.63611190184405e-14
+ pdiblcb = -0.025
+ drout = -2.03835735853155 ldrout = 1.66260803983147e-06 wdrout = 1.66443328246308e-06 pdrout = -1.12300195007201e-12
+ pscbe1 = 234237890.351731 lpscbe1 = 0.307796913526545 wpscbe1 = 29.6511740647848 ppscbe1 = -2.07900194053637e-7
+ pscbe2 = 1.17729860389986e-08 lpscbe2 = 2.01739268644305e-15 wpscbe2 = 1.85138462618454e-15 ppscbe2 = -1.36263982048721e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.76350543459814e-05 lalpha0 = 4.79702332198873e-11 walpha0 = 4.56838944623757e-11 palpha0 = -3.240130214744e-17
+ alpha1 = 7.42070134821428e-10 lalpha1 = -4.55388243122098e-16 walpha1 = -4.33683704284594e-16 palpha1 = 3.07590167263849e-22
+ beta0 = -235.917931284017 lbeta0 = 0.000169452542763189 wbeta0 = 0.000161376161014064 pbeta0 = -1.14456042199225e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.44159603248918e-06 lagidl = -5.87660224868919e-12 wagidl = -4.35088267549236e-12 pagidl = 3.9693277270493e-18
+ bgidl = -992180950.639868 lbgidl = 866.014098886511 wbgidl = 1364.8608653859 pbgidl = -0.000584945759036497
+ cgidl = 24766.5282614482 lcgidl = -0.0216227445599235 wcgidl = -0.0160570185973221 pcgidl = 1.46049963220221e-8
+ egidl = 7.30756299921459 legidl = -5.62985915410727e-06 wegidl = -4.32142849243674e-06 pegidl = 3.80266584620514e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 0.139534676118651 lkt1 = -2.14333985836712e-07 wkt1 = -6.14643736499889e-07 pkt1 = 3.29241439137551e-13
+ kt2 = -0.019032
+ at = 229339.026964286 lat = -0.15556620487442 wat = -0.0867367408569188 pat = 6.15180334527697e-8
+ ute = -1.3434125 lute = -9.67328343749999e-8
+ ua1 = 5.524e-10
+ ub1 = -4.57245346428571e-18 wub1 = 6.6298636123793e-25
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.86 pmos
* DC IV MOS Parameters
+ lmin = 6e-07 lmax = 8.0e-07 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.345600083238225+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -2.84286735553988e-07 wvth0 = -2.35348405101049e-07 pvth0 = 1.15038336457864e-13
+ k1 = 0.57315661187618 lk1 = 2.47894806270226e-08 wk1 = -2.7655072221193e-08 pk1 = -3.50905264952504e-15
+ k2 = 0.0291050296470879 lk2 = 5.08102747550879e-10 wk2 = 6.19758296132856e-09 pk2 = -5.00053353805815e-16
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 134531.170295577 lvsat = -0.0478616473464371 wvsat = -0.0289900008448478 pvsat = 2.31581832373675e-8
+ ua = 7.91066440498004e-09 lua = -3.70002764031288e-15 wua = -2.11214709450135e-15 pua = 1.18145752543688e-21
+ ub = -1.12137909662958e-17 lub = 6.92828875306842e-24 wub = 4.22952731530404e-24 pub = -2.42378048127152e-30
+ uc = -1.39893300407136e-12 luc = 5.69418078651683e-19 wuc = -8.61596644591578e-19 puc = -4.43283500710283e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0146135247201412 lu0 = -1.91669622105965e-10 wu0 = 2.72437589049307e-09 pu0 = -8.62130598940115e-16
+ a0 = -0.207347301027521 la0 = 6.4545193495285e-07 wa0 = 5.1737808555866e-07 pa0 = -3.49398244933507e-13
+ keta = 0.250220191756393 lketa = -2.03606746129757e-07 wketa = -1.21321730589239e-07 pketa = 8.80743979293742e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = -2.63759873785583 lags = 2.20392406086459e-06 wags = 1.17691064665417e-06 pags = -8.52631263168248e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '0.162013812530353+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -1.3422413476158e-07 wvoff = -1.06301381990881e-07 pvoff = 5.21598685553632e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '10.3673134818646+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -4.32529059918944e-06 wnfactor = -3.26523491972116e-06 pnfactor = 1.72285716336238e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 6.57536563392857e-05 lcit = -3.45348865532813e-11 wcit = -2.90593122722452e-11 pcit = 1.72274173966582e-17
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.93379884945137 leta0 = 9.42507553228316e-07 weta0 = 1.3567576706331e-06 peta0 = -6.55188173488013e-13
+ etab = -0.166187245348266 letab = 1.10447935435576e-07 wetab = 1.01853229772891e-07 petab = -6.9306801180686e-14
+ dsub = -0.373468212660117 ldsub = 3.35474447847452e-07 wdsub = 5.0943008472096e-07 pdsub = -2.57632685048049e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.49841646511415 lpclm = -5.61096181811415e-08 wpclm = -3.04864565512767e-07 ppclm = 9.71569835242463e-14
+ pdiblc1 = 0.255403744084621 lpdiblc1 = 3.51743959257796e-07 wpdiblc1 = 1.05704390801647e-07 ppdiblc1 = -1.73044894166074e-13
+ pdiblc2 = -0.0314101311255173 lpdiblc2 = 1.92493299685986e-08 wpdiblc2 = 1.82623666896451e-08 ppdiblc2 = -9.93432117015519e-15
+ pdiblcb = -0.025
+ drout = -2.47060246773729 ldrout = 1.96917788353565e-06 wdrout = 9.70423454204159e-07 pdrout = -6.3077547937937e-13
+ pscbe1 = -240203514.278644 lpscbe1 = 336.80536314762 wpscbe1 = 140.523335117 ppscbe1 = -7.88439804203377e-5
+ pscbe2 = 1.25399295264151e-08 lpscbe2 = 1.47343801799291e-15 wpscbe2 = 1.39203714674332e-15 ppscbe2 = -1.03684762069354e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000139105122503964 lalpha0 = 9.86603790609363e-11 walpha0 = 3.50230663091112e-11 palpha0 = -2.48401097797371e-17
+ alpha1 = 3.54625e-10 lalpha1 = -1.8059278125e-16
+ beta0 = -131.260013154095 lbeta0 = 9.52239143295422e-05 wbeta0 = 1.07127914776877e-05 pbeta0 = -7.59804735555001e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.35548247113527e-06 lagidl = 3.19972568000645e-12 wagidl = 4.23911646107348e-12 pagidl = -2.12312916056002e-18
+ bgidl = -4194888246.26064 lbgidl = 3137.53424830554 wbgidl = 2303.23640972826 pbgidl = -0.00125048861386132
+ cgidl = -18337.2382697941 lcgidl = 0.00894860185236016 wcgidl = 0.013391003031637 pcgidl = -6.28101301831722e-9
+ egidl = -3.27482114499542 legidl = 1.87569680017369e-06 wegidl = 2.75143023847538e-06 pegidl = -1.21375920869429e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = 1.04877751512 lkt1 = -8.59214469398419e-07 wkt1 = -5.85374985285981e-07 pkt1 = 3.08482577339087e-13
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.47310154375 lute = -4.75088009531244e-09 wute = -2.42896262201738e-07 pute = 1.72274173966582e-13
+ ua1 = 5.534185e-10 lua1 = -7.2237112499977e-19
+ ub1 = -1.14545940977232e-17 lub1 = 4.88115824426555e-24 wub1 = 2.35111538354e-24 pub1 = -1.19730550906775e-30
+ uc1 = -5.518905167685e-10 luc1 = 3.13978249018059e-16 wuc1 = 1.75060194094036e-16 puc1 = -1.24161442661195e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.87 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 6e-07 wmin = 4.2e-07 wmax = 7.0e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 4.5375e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 1.2277e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre)
+ toxe = '1.175e-08+MC_MM_SWITCH*GAU*(1.175e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre)
+ vth0 = '-0.690031318454674+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0 = -1.08885129020013e-07 wvth0 = -1.25090437296832e-07 pvth0 = 5.88894663535667e-14
+ k1 = 0.827591155466809 lk1 = -1.04781310696505e-07 wk1 = -6.72369549256842e-08 pk1 = 1.66480211177369e-14
+ k2 = -0.0693941075387678 lk2 = 5.06687883594479e-08 wk2 = 1.78001085450632e-08 pk2 = -6.40863950732271e-15
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -47730.1097866783 lvsat = 0.0449549095354516 wvsat = 0.0423606781503248 pvsat = -1.31771500409242e-8
+ ua = -6.66406354576978e-10 lua = 6.67845643991538e-16 wua = -1.44832982702827e-15 pua = 8.4340858197621e-22
+ ub = 1.9512301539758e-18 lub = 2.24001747570101e-25 wub = 3.9609933466648e-24 pub = -2.28702955774198e-30
+ uc = 8.08078287234235e-12 luc = -4.258127231412e-18 wuc = -1.17767854626666e-18 puc = -2.82318792282247e-25
+ rdsw = 788.47
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0104895406796788 lu0 = 1.9084692504995e-09 wu0 = 2.61153032819063e-09 pu0 = -8.04663996337597e-16
+ a0 = -1.20302893458061 la0 = 1.15250280683976e-06 wa0 = 1.71342329374369e-06 pa0 = -9.58484267201732e-13
+ keta = -0.34016648876305 lketa = 9.70476709247695e-08 wketa = 1.10267524552287e-07 pketa = -2.98624302514478e-14
+ a1 = 0.0
+ a2 = 0.5
+ ags = -1.01617130966482 lags = 1.37821214305832e-06 wags = 1.23377789891782e-06 pags = -8.81590911383512e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre)
+ voff = '-0.00825819193925859+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' lvoff = -4.75131164854306e-08 wvoff = -8.90874386687541e-08 pvoff = 4.33936679185699e-14
*(mismatch parameter sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre)
+ nfactor = '3.31169865068096+MC_MM_SWITCH*GAU*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor = -7.32218746409164e-07 wnfactor = -2.68930402526362e-07 pnfactor = 1.96989087980935e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -5.1423370625e-05 lcit = 2.51375144282813e-11 wcit = 2.42896262201738e-11 pcit = -9.94052953060611e-18
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = -1.07137221781493 leta0 = 5.03316791067456e-07 weta0 = 6.06971089862151e-07 peta0 = -2.73359357230406e-13
+ etab = 0.177976056575859 letab = -6.48172260692852e-08 wetab = -1.08127029466251e-07 petab = 3.76256458368471e-14
+ dsub = 0.408476767069836 ldsub = -6.27310330800269e-08 wdsub = -2.2070021383611e-08 pdsub = 1.30337439857038e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.12299661683596 lpclm = -8.83427060445474e-07 wpclm = -7.87864330413184e-07 ppclm = 3.43124613799784e-13
+ pdiblc1 = 5.28230638979032 lpdiblc1 = -2.20820621306783e-06 wpdiblc1 = -2.00450533301566e-06 ppdiblc1 = 9.01579407687891e-13
+ pdiblc2 = 0.0362915903430902 lpdiblc2 = -1.52277716892897e-08 wpdiblc2 = -1.91201190509867e-08 ppdiblc2 = 9.10270969326154e-15
+ pdiblcb = -0.025
+ drout = 2.0153149999156 ldrout = -3.1527558686659e-07 wdrout = -6.88792254866395e-07 pdrout = 2.1418012046481e-13
+ pscbe1 = 289922781.035108 lpscbe1 = 66.8385472590919 wpscbe1 = 74.3512172409605 ppscbe1 = -4.51458293919644e-5
+ pscbe2 = 1.8026849855846e-08 lpscbe2 = -1.32077615976978e-15 wpscbe2 = -3.11883498569308e-15 ppscbe2 = 1.26031401274971e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00014978930646844 lalpha0 = -4.84591088932604e-11 walpha0 = -3.70316908370358e-11 palpha0 = 1.18537752969382e-17
+ alpha1 = 0.0
+ beta0 = 74.5449543620496 lbeta0 = -9.5822653780546e-06 wbeta0 = -8.9606527784816e-06 pbeta0 = 2.42065413190422e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.01071367775527e-07 lagidl = 3.20216825620506e-13 wagidl = 3.80957249171881e-13 pagidl = -1.58361581899133e-19
+ bgidl = 2056754646.59452 lbgidl = -46.1148948809478 wbgidl = -333.72327666618 pbgidl = 9.23831064350506e-5
+ cgidl = -7750.50678138839 lcgidl = 0.00355730884188954 wcgidl = 0.00566483509326166 pcgidl = -2.34646199569957e-9
+ egidl = -0.432008666666309 legidl = 4.27994545584585e-07 wegidl = 1.00199839648804e-06 pegidl = -3.22861043162234e-13
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = -0.689872370390193 lkt1 = 2.61929847976478e-08 wkt1 = 3.29290201667861e-07 pkt1 = -1.57310669117157e-13
+ kt2 = -0.019032
+ at = 105600.770767857 lat = -0.0486846925135312 wat = -0.050751844437066 pat = 2.58453767795759e-8
+ ute = -1.90257537022857 lute = 2.13958666038901e-07 wute = 4.57683810561407e-07 pute = -1.8449622808805e-13
+ ua1 = 5.52e-10
+ ub1 = 1.94274678650001e-19 lub1 = -1.05102818010251e-24 wub1 = 8.41699820048573e-25 pub1 = -4.28635633359736e-31
+ uc1 = 1.167501147696e-09 luc1 = -5.61621956110488e-16 wuc1 = -6.14435994016312e-16 puc1 = 2.77889491134e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+40
+ noib = 8.5300000000000003e+24
+ noic = 84000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = 1.94170991e-10
+ cgso = 1.94170991e-10
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.8259105e-12
+ cgdl = 9.8259105e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 4.4983e-8
+ dwc = 0.0
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.00077934735
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = 9.9605453e-11
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = 1.47314e-10
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = '0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_g5v0d10v5
