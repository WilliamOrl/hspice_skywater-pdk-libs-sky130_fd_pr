* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* ./models_capacitors.spice created from ./models.spice
*

.param GAU = AGAUSS(0,1.0,1)

**********************************
******************************************************************
******************************************************************
********************************************************************
*          model for interconnect capacitance                      *
********************************************************************

***************************************
** minimum width for different layers *
***************************************

.param
+ wminp1= 0.15u
+ wminl1= 0.14u
+ wminm1= 0.14u
+ wminm2= 0.14u
+ wminm3= 0.3u
+ wminm4= 0.3u
+ wminm5= 0.8u
+ wminrdl= 10.0u

.model mcp1f c tc1 = 0 tc2 = 0 cox = 'cp1f' capsw = 'cp1fsw' w = 'wminp1' tref = 25

.model mcl1f c tc1 = 0 tc2 = 0 cox = 'cl1f' capsw = 'cl1fsw' w = 'wminl1' tref = 25
.model mcl1d c tc1 = 0 tc2 = 0 cox = 'cl1d' capsw = 'cl1dsw' w = 'wminl1' tref = 25
.model mcl1p1 c tc1 = 0 tc2 = 0 cox = 'cl1p1' capsw = 'cl1p1sw' w = 'wminl1' tref = 25

.model mcm1f c tc1 = 0 tc2 = 0 cox = 'cm1f' capsw = 'cm1fsw' w = 'wminm1' tref = 25
.model mcm1d c tc1 = 0 tc2 = 0 cox = 'cm1d' capsw = 'cm1dsw' w = 'wminm1' tref = 25
.model mcm1p1 c tc1 = 0 tc2 = 0 cox = 'cm1p1' capsw = 'cm1p1sw' w = 'wminm1' tref = 25
.model mcm1l1 c tc1 = 0 tc2 = 0 cox = 'cm1l1' capsw = 'cm1l1sw' w = 'wminm1' tref = 25

.model mcm2f c tc1 = 0 tc2 = 0 cox = 'cm2f' capsw = 'cm2fsw' w = 'wminm2' tref = 25
.model mcm2d c tc1 = 0 tc2 = 0 cox = 'cm2d' capsw = 'cm2dsw' w = 'wminm2' tref = 25
.model mcm2p1 c tc1 = 0 tc2 = 0 cox = 'cm2p1' capsw = 'cm2p1sw' w = 'wminm2' tref = 25
.model mcm2l1 c tc1 = 0 tc2 = 0 cox = 'cm2l1' capsw = 'cm2l1sw' w = 'wminm2' tref = 25
.model mcm2m1 c tc1 = 0 tc2 = 0 cox = 'cm2m1' capsw = 'cm2m1sw' w = 'wminm2' tref = 25

.model mcm3f c tc1 = 0 tc2 = 0 cox = 'cm3f' capsw = 'cm3fsw' w = 'wminm3' tref = 25
.model mcm3d c tc1 = 0 tc2 = 0 cox = 'cm3d' capsw = 'cm3dsw' w = 'wminm3' tref = 25
.model mcm3p1 c tc1 = 0 tc2 = 0 cox = 'cm3p1' capsw = 'cm3p1sw' w = 'wminm3' tref = 25
.model mcm3l1 c tc1 = 0 tc2 = 0 cox = 'cm3l1' capsw = 'cm3l1sw' w = 'wminm3' tref = 25
.model mcm3m1 c tc1 = 0 tc2 = 0 cox = 'cm3m1' capsw = 'cm3m1sw' w = 'wminm3' tref = 25
.model mcm3m2 c tc1 = 0 tc2 = 0 cox = 'cm3m2' capsw = 'cm3m2sw' w = 'wminm3' tref = 25

.model mcm4f c tc1 = 0 tc2 = 0 cox = 'cm4f' capsw = 'cm4fsw' w = 'wminm4' tref = 25
.model mcm4d c tc1 = 0 tc2 = 0 cox = 'cm4d' capsw = 'cm4dsw' w = 'wminm4' tref = 25
.model mcm4p1 c tc1 = 0 tc2 = 0 cox = 'cm4p1' capsw = 'cm4p1sw' w = 'wminm4' tref = 25
.model mcm4l1 c tc1 = 0 tc2 = 0 cox = 'cm4l1' capsw = 'cm4l1sw' w = 'wminm4' tref = 25
.model mcm4m1 c tc1 = 0 tc2 = 0 cox = 'cm4m1' capsw = 'cm4m1sw' w = 'wminm4' tref = 25
.model mcm4m2 c tc1 = 0 tc2 = 0 cox = 'cm4m2' capsw = 'cm4m2sw' w = 'wminm4' tref = 25
.model mcm4m3 c tc1 = 0 tc2 = 0 cox = 'cm4m3' capsw = 'cm4m3sw' w = 'wminm4' tref = 25

.model mcm5f c tc1 = 0 tc2 = 0 cox = 'cm5f' capsw = 'cm5fsw' w = 'wminm5' tref = 25
.model mcm5d c tc1 = 0 tc2 = 0 cox = 'cm5d' capsw = 'cm5dsw' w = 'wminm5' tref = 25
.model mcm5p1 c tc1 = 0 tc2 = 0 cox = 'cm5p1' capsw = 'cm5p1sw' w = 'wminm5' tref = 25
.model mcm5l1 c tc1 = 0 tc2 = 0 cox = 'cm5l1' capsw = 'cm5l1sw' w = 'wminm5' tref = 25
.model mcm5m1 c tc1 = 0 tc2 = 0 cox = 'cm5m1' capsw = 'cm5m1sw' w = 'wminm5' tref = 25
.model mcm5m2 c tc1 = 0 tc2 = 0 cox = 'cm5m2' capsw = 'cm5m2sw' w = 'wminm5' tref = 25
.model mcm5m3 c tc1 = 0 tc2 = 0 cox = 'cm5m3' capsw = 'cm5m3sw' w = 'wminm5' tref = 25
.model mcm5m4 c tc1 = 0 tc2 = 0 cox = 'cm5m4' capsw = 'cm5m4sw' w = 'wminm5' tref = 25

.model mcrdlf c tc1 = 0 tc2 = 0 cox = 'crdlf' capsw = 'crdlfsw' w = 'wminrdl' tref = 25
.model mcrdld c tc1 = 0 tc2 = 0 cox = 'crdld' capsw = 'crdldsw' w = 'wminrdl' tref = 25
.model mcrdlp1 c tc1 = 0 tc2 = 0 cox = 'crdlp1' capsw = 'crdlp1sw' w = 'wminrdl' tref = 25
.model mcrdll1 c tc1 = 0 tc2 = 0 cox = 'crdll1' capsw = 'crdll1sw' w = 'wminrdl' tref = 25
.model mcrdlm1 c tc1 = 0 tc2 = 0 cox = 'crdlm1' capsw = 'crdlm1sw' w = 'wminrdl' tref = 25
.model mcrdlm2 c tc1 = 0 tc2 = 0 cox = 'crdlm2' capsw = 'crdlm2sw' w = 'wminrdl' tref = 25
.model mcrdlm3 c tc1 = 0 tc2 = 0 cox = 'crdlm3' capsw = 'crdlm3sw' w = 'wminrdl' tref = 25
.model mcrdlm4 c tc1 = 0 tc2 = 0 cox = 'crdlm4' capsw = 'crdlm4sw' w = 'wminrdl' tref = 25
.model mcrdlm5 c tc1 = 0 tc2 = 0 cox = 'crdlm5' capsw = 'crdlm5sw' w = 'wminrdl' tref = 25

******************************************************************
******************************************************************
*  *****************************************************
*  12/03/2020 Usman Suriono
*      Why     : New model structure
*      What    : Converted from MIMCap models
*
*  *****************************************************
*
*  MIM Capacitor Model
*  -----------------------------------------------------

.subckt  sky130_fd_pr__cap_mim_m3_1 c0 c1  mult=1
+ w=1 l=1
+ 
.param  wc = 'w+sw_cap_mim_dw*1e6'
+ lc = 'l+sw_cap_mim_dw*1e6'
+ carea = 'sw_cap_mim_ca*wc*lc*(1+mismatch_factor*MC_MM_SWITCH*GAU*sw_mm_cmim/sqrt(wc*lc*mult))'

c1 c0  c1 c = 'carea'


.ends sky130_fd_pr__cap_mim_m3_1

*  -----------------------------------------------------

.subckt  sky130_fd_pr__cap_mim_m3_2 c0 c1  mult=1
+ w=1 l=1
+ 
.param  wc = 'w+sw_cap_mim_dw*1e6'
+ lc = 'l+sw_cap_mim_dw*1e6'
+ carea = 'sw_cap_mim_ca*wc*lc*(1+mismatch_factor*MC_MM_SWITCH*GAU*sw_mm_cmim/sqrt(wc*lc*mult))'

c1 c0  c1 c = 'carea'


.ends sky130_fd_pr__cap_mim_m3_2

******************************************************************
******************************************************************
* *************************** Poly Resistor Parasitic Capacitance to Substrate ************************
* 2021/02/14  UZMN (Usman Suriono)
*      Why  : New parasitic capacitance from Poly to silicon over thick STI oxide
*      What : Copied from but changed the cap/area from 1.53e-4 to 1.06e-4
*             Poly resistors sit on STI with the thickness of 3262A, i.e 1.06e-4 F/m^2

.subckt  sky130_fd_pr__model__parasitic__cap_p2ps r0 sub mult=1
+ w=1 l=1
+ 
.param  crpf_precision = 1.06e-04

c0 r0 sub  c = 'l*w*crpf_precision*1e-12*sw_fox_poly_cap'


.ends sky130_fd_pr__model__parasitic__cap_p2ps
